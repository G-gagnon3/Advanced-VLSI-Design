
module FIR (input logic clk, reset, input logic [31:0] val_in, output logic [31:0] val_out);
  logic [3199:0] history;
  logic [6511:0] value_grid;
  logic [31:0] cur_val_q;
  logic [12831:0] tap_outputs;
  logic [31:0] val_out_buffer;
  assign value_grid = {history, cur_val_q};
  assign cur_val_q = val_in;
  always_comb begin
    logic [6415:0] adder_tree_tier_0_p0_in;
    logic [3215:0] adder_tree_tier_1_p0_in;
    logic [1615:0] adder_tree_tier_2_p0_in;
    logic [815:0] adder_tree_tier_3_p0_in;
    logic [415:0] adder_tree_tier_4_p0_in;
    logic [207:0] adder_tree_tier_5_p0_in;
    logic [111:0] adder_tree_tier_6_p0_in;
    logic [63:0] adder_tree_tier_7_p0_in;
    logic [31:0] adder_tree_tier_8_p0_in;
    logic [15:0] adder_tree_tier_9_p0_in;
    logic [6415:0] adder_tree_tier_0_p1_in;
    logic [3215:0] adder_tree_tier_1_p1_in;
    logic [1615:0] adder_tree_tier_2_p1_in;
    logic [815:0] adder_tree_tier_3_p1_in;
    logic [415:0] adder_tree_tier_4_p1_in;
    logic [207:0] adder_tree_tier_5_p1_in;
    logic [111:0] adder_tree_tier_6_p1_in;
    logic [63:0] adder_tree_tier_7_p1_in;
    logic [31:0] adder_tree_tier_8_p1_in;
    logic [15:0] adder_tree_tier_9_p1_in;
    tap_outputs[15:0] = value_grid[47:32] * 11390;
    tap_outputs[31:16] = value_grid[63:48] * 11392;
    tap_outputs[6463:6448] = value_grid[79:64] * 11391;
    tap_outputs[6479:6464] = value_grid[95:80] * 11391;
    tap_outputs[6495:6480] = value_grid[111:96] * 11391;
    tap_outputs[95:80] = value_grid[127:112] * 11390;
    tap_outputs[6527:6512] = value_grid[143:128] * 11389;
    tap_outputs[6543:6528] = value_grid[159:144] * 11389;
    tap_outputs[6559:6544] = value_grid[175:160] * 11389;
    tap_outputs[159:144] = value_grid[191:176] * 11390;
    tap_outputs[6591:6576] = value_grid[207:192] * 11391;
    tap_outputs[191:176] = value_grid[223:208] * 11392;
    tap_outputs[6623:6608] = value_grid[239:224] * 11393;
    tap_outputs[223:208] = value_grid[255:240] * 11392;
    tap_outputs[239:224] = value_grid[271:256] * 11390;
    tap_outputs[255:240] = value_grid[287:272] * 11388;
    tap_outputs[6687:6672] = value_grid[303:288] * 11387;
    tap_outputs[6703:6688] = value_grid[319:304] * 11387;
    tap_outputs[6719:6704] = value_grid[335:320] * 11389;
    tap_outputs[319:304] = value_grid[351:336] * 11392;
    tap_outputs[335:320] = value_grid[367:352] * 11394;
    tap_outputs[351:336] = value_grid[383:368] * 11396;
    tap_outputs[6783:6768] = value_grid[399:384] * 11395;
    tap_outputs[6799:6784] = value_grid[415:400] * 11391;
    tap_outputs[6815:6800] = value_grid[431:416] * 11387;
    tap_outputs[415:400] = value_grid[447:432] * 11384;
    tap_outputs[6847:6832] = value_grid[463:448] * 11383;
    tap_outputs[447:432] = value_grid[479:464] * 11386;
    tap_outputs[6879:6864] = value_grid[495:480] * 11391;
    tap_outputs[6895:6880] = value_grid[511:496] * 11397;
    tap_outputs[495:480] = value_grid[527:512] * 11400;
    tap_outputs[511:496] = value_grid[543:528] * 11400;
    tap_outputs[6943:6928] = value_grid[559:544] * 11395;
    tap_outputs[6959:6944] = value_grid[575:560] * 11387;
    tap_outputs[559:544] = value_grid[591:576] * 11380;
    tap_outputs[6991:6976] = value_grid[607:592] * 11377;
    tap_outputs[591:576] = value_grid[623:608] * 11380;
    tap_outputs[607:592] = value_grid[639:624] * 11388;
    tap_outputs[7039:7024] = value_grid[655:640] * 11399;
    tap_outputs[7055:7040] = value_grid[671:656] * 11407;
    tap_outputs[655:640] = value_grid[687:672] * 11408;
    tap_outputs[7087:7072] = value_grid[703:688] * 11401;
    tap_outputs[687:672] = value_grid[719:704] * 11388;
    tap_outputs[7119:7104] = value_grid[735:720] * 11375;
    tap_outputs[7135:7120] = value_grid[751:736] * 11367;
    tap_outputs[7151:7136] = value_grid[767:752] * 11369;
    tap_outputs[7167:7152] = value_grid[783:768] * 11381;
    tap_outputs[7183:7168] = value_grid[799:784] * 11399;
    tap_outputs[7199:7184] = value_grid[815:800] * 11415;
    tap_outputs[7215:7200] = value_grid[831:816] * 11421;
    tap_outputs[7231:7216] = value_grid[847:832] * 11413;
    tap_outputs[831:816] = value_grid[863:848] * 11394;
    tap_outputs[7263:7248] = value_grid[879:864] * 11371;
    tap_outputs[7279:7264] = value_grid[895:880] * 11355;
    tap_outputs[7295:7280] = value_grid[911:896] * 11353;
    tap_outputs[7311:7296] = value_grid[927:912] * 11369;
    tap_outputs[911:896] = value_grid[943:928] * 11396;
    tap_outputs[7343:7328] = value_grid[959:944] * 11423;
    tap_outputs[943:928] = value_grid[975:960] * 11438;
    tap_outputs[7375:7360] = value_grid[991:976] * 11433;
    tap_outputs[7391:7376] = value_grid[1007:992] * 11407;
    tap_outputs[7407:7392] = value_grid[1023:1008] * 11371;
    tap_outputs[7423:7408] = value_grid[1039:1024] * 11341;
    tap_outputs[1023:1008] = value_grid[1055:1040] * 11330;
    tap_outputs[7455:7440] = value_grid[1071:1056] * 11347;
    tap_outputs[7471:7456] = value_grid[1087:1072] * 11385;
    tap_outputs[7487:7472] = value_grid[1103:1088] * 11429;
    tap_outputs[1087:1072] = value_grid[1119:1104] * 11460;
    tap_outputs[7519:7504] = value_grid[1135:1120] * 11461;
    tap_outputs[1119:1104] = value_grid[1151:1136] * 11430;
    tap_outputs[1135:1120] = value_grid[1167:1152] * 11378;
    tap_outputs[7567:7552] = value_grid[1183:1168] * 11327;
    tap_outputs[7583:7568] = value_grid[1199:1184] * 11301;
    tap_outputs[1183:1168] = value_grid[1215:1200] * 11314;
    tap_outputs[7615:7600] = value_grid[1231:1216] * 11363;
    tap_outputs[7631:7616] = value_grid[1247:1232] * 11429;
    tap_outputs[7647:7632] = value_grid[1263:1248] * 11483;
    tap_outputs[7663:7648] = value_grid[1279:1264] * 11499;
    tap_outputs[7679:7664] = value_grid[1295:1280] * 11467;
    tap_outputs[1279:1264] = value_grid[1311:1296] * 11396;
    tap_outputs[7711:7696] = value_grid[1327:1312] * 11317;
    tap_outputs[1311:1296] = value_grid[1343:1328] * 11266;
    tap_outputs[7743:7728] = value_grid[1359:1344] * 11267;
    tap_outputs[7759:7744] = value_grid[1375:1360] * 11325;
    tap_outputs[7775:7760] = value_grid[1391:1376] * 11417;
    tap_outputs[7791:7776] = value_grid[1407:1392] * 11505;
    tap_outputs[7807:7792] = value_grid[1423:1408] * 11547;
    tap_outputs[7823:7808] = value_grid[1439:1424] * 11521;
    tap_outputs[7839:7824] = value_grid[1455:1440] * 11433;
    tap_outputs[7855:7840] = value_grid[1471:1456] * 11319;
    tap_outputs[7871:7856] = value_grid[1487:1472] * 11229;
    tap_outputs[1471:1456] = value_grid[1503:1488] * 11206;
    tap_outputs[1487:1472] = value_grid[1519:1504] * 11266;
    tap_outputs[7919:7904] = value_grid[1535:1520] * 11387;
    tap_outputs[7935:7920] = value_grid[1551:1536] * 11519;
    tap_outputs[1535:1520] = value_grid[1567:1552] * 11602;
    tap_outputs[1551:1536] = value_grid[1583:1568] * 11594;
    tap_outputs[7983:7968] = value_grid[1599:1584] * 11493;
    tap_outputs[1583:1568] = value_grid[1615:1600] * 11338;
    tap_outputs[1599:1584] = value_grid[1631:1616] * 11196;
    tap_outputs[1615:1600] = value_grid[1647:1632] * 11132;
    tap_outputs[8047:8032] = value_grid[1663:1648] * 11181;
    tap_outputs[1647:1632] = value_grid[1679:1664] * 11330;
    tap_outputs[1663:1648] = value_grid[1695:1680] * 11516;
    tap_outputs[1679:1664] = value_grid[1711:1696] * 11658;
    tap_outputs[1695:1680] = value_grid[1727:1712] * 11688;
    tap_outputs[1711:1696] = value_grid[1743:1728] * 11584;
    tap_outputs[1727:1712] = value_grid[1759:1744] * 11386;
    tap_outputs[1743:1728] = value_grid[1775:1760] * 11176;
    tap_outputs[8175:8160] = value_grid[1791:1776] * 11049;
    tap_outputs[8191:8176] = value_grid[1807:1792] * 11069;
    tap_outputs[8207:8192] = value_grid[1823:1808] * 11237;
    tap_outputs[8223:8208] = value_grid[1839:1824] * 11485;
    tap_outputs[8239:8224] = value_grid[1855:1840] * 11707;
    tap_outputs[8255:8240] = value_grid[1871:1856] * 11799;
    tap_outputs[1855:1840] = value_grid[1887:1872] * 11712;
    tap_outputs[8287:8272] = value_grid[1903:1888] * 11473;
    tap_outputs[1887:1872] = value_grid[1919:1904] * 11180;
    tap_outputs[8319:8304] = value_grid[1935:1920] * 10965;
    tap_outputs[8335:8320] = value_grid[1951:1936] * 10929;
    tap_outputs[1935:1920] = value_grid[1967:1952] * 11100;
    tap_outputs[1951:1936] = value_grid[1983:1968] * 11414;
    tap_outputs[8383:8368] = value_grid[1999:1984] * 11737;
    tap_outputs[1983:1968] = value_grid[2015:2000] * 11924;
    tap_outputs[1999:1984] = value_grid[2031:2016] * 11880;
    tap_outputs[8431:8416] = value_grid[2047:2032] * 11611;
    tap_outputs[8447:8432] = value_grid[2063:2048] * 11225;
    tap_outputs[8463:8448] = value_grid[2079:2064] * 10891;
    tap_outputs[8479:8464] = value_grid[2095:2080] * 10761;
    tap_outputs[2079:2064] = value_grid[2111:2096] * 10910;
    tap_outputs[8511:8496] = value_grid[2127:2112] * 11285;
    tap_outputs[8527:8512] = value_grid[2143:2128] * 11731;
    tap_outputs[8543:8528] = value_grid[2159:2144] * 12051;
    tap_outputs[2143:2128] = value_grid[2175:2160] * 12090;
    tap_outputs[8575:8560] = value_grid[2191:2176] * 11815;
    tap_outputs[2175:2160] = value_grid[2207:2192] * 11330;
    tap_outputs[2191:2176] = value_grid[2223:2208] * 10842;
    tap_outputs[8623:8608] = value_grid[2239:2224] * 10573;
    tap_outputs[2223:2208] = value_grid[2255:2240] * 10658;
    tap_outputs[2239:2224] = value_grid[2271:2256] * 11080;
    tap_outputs[8671:8656] = value_grid[2287:2272] * 11669;
    tap_outputs[2271:2256] = value_grid[2303:2288] * 12168;
    tap_outputs[8703:8688] = value_grid[2319:2304] * 12345;
    tap_outputs[8719:8704] = value_grid[2335:2320] * 12101;
    tap_outputs[8735:8720] = value_grid[2351:2336] * 11519;
    tap_outputs[2335:2320] = value_grid[2367:2352] * 10842;
    tap_outputs[2351:2336] = value_grid[2383:2368] * 10372;
    tap_outputs[2367:2352] = value_grid[2399:2384] * 10334;
    tap_outputs[8799:8784] = value_grid[2415:2400] * 10773;
    tap_outputs[2399:2384] = value_grid[2431:2416] * 11520;
    tap_outputs[8831:8816] = value_grid[2447:2432] * 12255;
    tap_outputs[8847:8832] = value_grid[2463:2448] * 12645;
    tap_outputs[2447:2432] = value_grid[2479:2464] * 12490;
    tap_outputs[2463:2448] = value_grid[2495:2480] * 11826;
    tap_outputs[8895:8880] = value_grid[2511:2496] * 10921;
    tap_outputs[2495:2480] = value_grid[2527:2512] * 10170;
    tap_outputs[8927:8912] = value_grid[2543:2528] * 9923;
    tap_outputs[8943:8928] = value_grid[2559:2544] * 10327;
    tap_outputs[8959:8944] = value_grid[2575:2560] * 11241;
    tap_outputs[8975:8960] = value_grid[2591:2576] * 12285;
    tap_outputs[8991:8976] = value_grid[2607:2592] * 12995;
    tap_outputs[9007:8992] = value_grid[2623:2608] * 13023;
    tap_outputs[9023:9008] = value_grid[2639:2624] * 12311;
    tap_outputs[2623:2608] = value_grid[2655:2640] * 11128;
    tap_outputs[9055:9040] = value_grid[2671:2656] * 9979;
    tap_outputs[2655:2640] = value_grid[2687:2672] * 9388;
    tap_outputs[9087:9072] = value_grid[2703:2688] * 9667;
    tap_outputs[2687:2672] = value_grid[2719:2704] * 10754;
    tap_outputs[2703:2688] = value_grid[2735:2720] * 12216;
    tap_outputs[2719:2704] = value_grid[2751:2736] * 13416;
    tap_outputs[9151:9136] = value_grid[2767:2752] * 13787;
    tap_outputs[9167:9152] = value_grid[2783:2768] * 13091;
    tap_outputs[9183:9168] = value_grid[2799:2784] * 11557;
    tap_outputs[2783:2768] = value_grid[2815:2800] * 9812;
    tap_outputs[9215:9200] = value_grid[2831:2816] * 8637;
    tap_outputs[9231:9216] = value_grid[2847:2832] * 8619;
    tap_outputs[9247:9232] = value_grid[2863:2848] * 9877;
    tap_outputs[2847:2832] = value_grid[2879:2864] * 11956;
    tap_outputs[9279:9264] = value_grid[2895:2880] * 13985;
    tap_outputs[2879:2864] = value_grid[2911:2896] * 15028;
    tap_outputs[2895:2880] = value_grid[2927:2912] * 14498;
    tap_outputs[9327:9312] = value_grid[2943:2928] * 12463;
    tap_outputs[9343:9328] = value_grid[2959:2944] * 9683;
    tap_outputs[2943:2928] = value_grid[2975:2960] * 7350;
    tap_outputs[2959:2944] = value_grid[2991:2976] * 6602;
    tap_outputs[9391:9376] = value_grid[3007:2992] * 8001;
    tap_outputs[9407:9392] = value_grid[3023:3008] * 11213;
    tap_outputs[3007:2992] = value_grid[3039:3024] * 15026;
    tap_outputs[3023:3008] = value_grid[3055:3040] * 17762;
    tap_outputs[9455:9440] = value_grid[3071:3056] * 17947;
    tap_outputs[3055:3040] = value_grid[3087:3072] * 14992;
    tap_outputs[9487:9472] = value_grid[3103:3088] * 9601;
    tap_outputs[9503:9488] = value_grid[3119:3104] * 3723;
    tap_outputs[3103:3088] = value_grid[3135:3120] * 0;
    tap_outputs[3119:3104] = value_grid[3151:3136] * 874;
    tap_outputs[9551:9536] = value_grid[3167:3152] * 7657;
    tap_outputs[9567:9552] = value_grid[3183:3168] * 19907;
    tap_outputs[3167:3152] = value_grid[3199:3184] * 35362;
    tap_outputs[9599:9584] = value_grid[3215:3200] * 50489;
    tap_outputs[9615:9600] = value_grid[3231:3216] * 61505;
    tap_outputs[9631:9616] = value_grid[3247:3232] * 65535;
    tap_outputs[9647:9632] = value_grid[3263:3248] * 61505;
    tap_outputs[9663:9648] = value_grid[3279:3264] * 50489;
    tap_outputs[3263:3248] = value_grid[3295:3280] * 35362;
    tap_outputs[9695:9680] = value_grid[3311:3296] * 19907;
    tap_outputs[9711:9696] = value_grid[3327:3312] * 7657;
    tap_outputs[3311:3296] = value_grid[3343:3328] * 874;
    tap_outputs[3327:3312] = value_grid[3359:3344] * 0;
    tap_outputs[9759:9744] = value_grid[3375:3360] * 3723;
    tap_outputs[9775:9760] = value_grid[3391:3376] * 9601;
    tap_outputs[3375:3360] = value_grid[3407:3392] * 14992;
    tap_outputs[9807:9792] = value_grid[3423:3408] * 17947;
    tap_outputs[3407:3392] = value_grid[3439:3424] * 17762;
    tap_outputs[3423:3408] = value_grid[3455:3440] * 15026;
    tap_outputs[9855:9840] = value_grid[3471:3456] * 11213;
    tap_outputs[9871:9856] = value_grid[3487:3472] * 8001;
    tap_outputs[3471:3456] = value_grid[3503:3488] * 6602;
    tap_outputs[3487:3472] = value_grid[3519:3504] * 7350;
    tap_outputs[9919:9904] = value_grid[3535:3520] * 9683;
    tap_outputs[9935:9920] = value_grid[3551:3536] * 12463;
    tap_outputs[3535:3520] = value_grid[3567:3552] * 14498;
    tap_outputs[3551:3536] = value_grid[3583:3568] * 15028;
    tap_outputs[9983:9968] = value_grid[3599:3584] * 13985;
    tap_outputs[3583:3568] = value_grid[3615:3600] * 11956;
    tap_outputs[10015:10000] = value_grid[3631:3616] * 9877;
    tap_outputs[10031:10016] = value_grid[3647:3632] * 8619;
    tap_outputs[10047:10032] = value_grid[3663:3648] * 8637;
    tap_outputs[3647:3632] = value_grid[3679:3664] * 9812;
    tap_outputs[10079:10064] = value_grid[3695:3680] * 11557;
    tap_outputs[10095:10080] = value_grid[3711:3696] * 13091;
    tap_outputs[10111:10096] = value_grid[3727:3712] * 13787;
    tap_outputs[3711:3696] = value_grid[3743:3728] * 13416;
    tap_outputs[3727:3712] = value_grid[3759:3744] * 12216;
    tap_outputs[3743:3728] = value_grid[3775:3760] * 10754;
    tap_outputs[10175:10160] = value_grid[3791:3776] * 9667;
    tap_outputs[3775:3760] = value_grid[3807:3792] * 9388;
    tap_outputs[10207:10192] = value_grid[3823:3808] * 9979;
    tap_outputs[3807:3792] = value_grid[3839:3824] * 11128;
    tap_outputs[10239:10224] = value_grid[3855:3840] * 12311;
    tap_outputs[10255:10240] = value_grid[3871:3856] * 13023;
    tap_outputs[10271:10256] = value_grid[3887:3872] * 12995;
    tap_outputs[10287:10272] = value_grid[3903:3888] * 12285;
    tap_outputs[10303:10288] = value_grid[3919:3904] * 11241;
    tap_outputs[10319:10304] = value_grid[3935:3920] * 10327;
    tap_outputs[10335:10320] = value_grid[3951:3936] * 9923;
    tap_outputs[3935:3920] = value_grid[3967:3952] * 10170;
    tap_outputs[10367:10352] = value_grid[3983:3968] * 10921;
    tap_outputs[3967:3952] = value_grid[3999:3984] * 11826;
    tap_outputs[3983:3968] = value_grid[4015:4000] * 12490;
    tap_outputs[10415:10400] = value_grid[4031:4016] * 12645;
    tap_outputs[10431:10416] = value_grid[4047:4032] * 12255;
    tap_outputs[4031:4016] = value_grid[4063:4048] * 11520;
    tap_outputs[10463:10448] = value_grid[4079:4064] * 10773;
    tap_outputs[4063:4048] = value_grid[4095:4080] * 10334;
    tap_outputs[4079:4064] = value_grid[4111:4096] * 10372;
    tap_outputs[4095:4080] = value_grid[4127:4112] * 10842;
    tap_outputs[10527:10512] = value_grid[4143:4128] * 11519;
    tap_outputs[10543:10528] = value_grid[4159:4144] * 12101;
    tap_outputs[10559:10544] = value_grid[4175:4160] * 12345;
    tap_outputs[4159:4144] = value_grid[4191:4176] * 12168;
    tap_outputs[10591:10576] = value_grid[4207:4192] * 11669;
    tap_outputs[4191:4176] = value_grid[4223:4208] * 11080;
    tap_outputs[4207:4192] = value_grid[4239:4224] * 10658;
    tap_outputs[10639:10624] = value_grid[4255:4240] * 10573;
    tap_outputs[4239:4224] = value_grid[4271:4256] * 10842;
    tap_outputs[4255:4240] = value_grid[4287:4272] * 11330;
    tap_outputs[10687:10672] = value_grid[4303:4288] * 11815;
    tap_outputs[4287:4272] = value_grid[4319:4304] * 12090;
    tap_outputs[10719:10704] = value_grid[4335:4320] * 12051;
    tap_outputs[10735:10720] = value_grid[4351:4336] * 11731;
    tap_outputs[10751:10736] = value_grid[4367:4352] * 11285;
    tap_outputs[4351:4336] = value_grid[4383:4368] * 10910;
    tap_outputs[10783:10768] = value_grid[4399:4384] * 10761;
    tap_outputs[10799:10784] = value_grid[4415:4400] * 10891;
    tap_outputs[10815:10800] = value_grid[4431:4416] * 11225;
    tap_outputs[10831:10816] = value_grid[4447:4432] * 11611;
    tap_outputs[4431:4416] = value_grid[4463:4448] * 11880;
    tap_outputs[4447:4432] = value_grid[4479:4464] * 11924;
    tap_outputs[10879:10864] = value_grid[4495:4480] * 11737;
    tap_outputs[4479:4464] = value_grid[4511:4496] * 11414;
    tap_outputs[4495:4480] = value_grid[4527:4512] * 11100;
    tap_outputs[10927:10912] = value_grid[4543:4528] * 10929;
    tap_outputs[10943:10928] = value_grid[4559:4544] * 10965;
    tap_outputs[4543:4528] = value_grid[4575:4560] * 11180;
    tap_outputs[10975:10960] = value_grid[4591:4576] * 11473;
    tap_outputs[4575:4560] = value_grid[4607:4592] * 11712;
    tap_outputs[11007:10992] = value_grid[4623:4608] * 11799;
    tap_outputs[11023:11008] = value_grid[4639:4624] * 11707;
    tap_outputs[11039:11024] = value_grid[4655:4640] * 11485;
    tap_outputs[11055:11040] = value_grid[4671:4656] * 11237;
    tap_outputs[11071:11056] = value_grid[4687:4672] * 11069;
    tap_outputs[11087:11072] = value_grid[4703:4688] * 11049;
    tap_outputs[4687:4672] = value_grid[4719:4704] * 11176;
    tap_outputs[4703:4688] = value_grid[4735:4720] * 11386;
    tap_outputs[4719:4704] = value_grid[4751:4736] * 11584;
    tap_outputs[4735:4720] = value_grid[4767:4752] * 11688;
    tap_outputs[4751:4736] = value_grid[4783:4768] * 11658;
    tap_outputs[4767:4752] = value_grid[4799:4784] * 11516;
    tap_outputs[4783:4768] = value_grid[4815:4800] * 11330;
    tap_outputs[11215:11200] = value_grid[4831:4816] * 11181;
    tap_outputs[4815:4800] = value_grid[4847:4832] * 11132;
    tap_outputs[4831:4816] = value_grid[4863:4848] * 11196;
    tap_outputs[4847:4832] = value_grid[4879:4864] * 11338;
    tap_outputs[11279:11264] = value_grid[4895:4880] * 11493;
    tap_outputs[4879:4864] = value_grid[4911:4896] * 11594;
    tap_outputs[4895:4880] = value_grid[4927:4912] * 11602;
    tap_outputs[11327:11312] = value_grid[4943:4928] * 11519;
    tap_outputs[11343:11328] = value_grid[4959:4944] * 11387;
    tap_outputs[4943:4928] = value_grid[4975:4960] * 11266;
    tap_outputs[4959:4944] = value_grid[4991:4976] * 11206;
    tap_outputs[11391:11376] = value_grid[5007:4992] * 11229;
    tap_outputs[11407:11392] = value_grid[5023:5008] * 11319;
    tap_outputs[11423:11408] = value_grid[5039:5024] * 11433;
    tap_outputs[11439:11424] = value_grid[5055:5040] * 11521;
    tap_outputs[11455:11440] = value_grid[5071:5056] * 11547;
    tap_outputs[11471:11456] = value_grid[5087:5072] * 11505;
    tap_outputs[11487:11472] = value_grid[5103:5088] * 11417;
    tap_outputs[11503:11488] = value_grid[5119:5104] * 11325;
    tap_outputs[11519:11504] = value_grid[5135:5120] * 11267;
    tap_outputs[5119:5104] = value_grid[5151:5136] * 11266;
    tap_outputs[11551:11536] = value_grid[5167:5152] * 11317;
    tap_outputs[5151:5136] = value_grid[5183:5168] * 11396;
    tap_outputs[11583:11568] = value_grid[5199:5184] * 11467;
    tap_outputs[11599:11584] = value_grid[5215:5200] * 11499;
    tap_outputs[11615:11600] = value_grid[5231:5216] * 11483;
    tap_outputs[11631:11616] = value_grid[5247:5232] * 11429;
    tap_outputs[11647:11632] = value_grid[5263:5248] * 11363;
    tap_outputs[5247:5232] = value_grid[5279:5264] * 11314;
    tap_outputs[11679:11664] = value_grid[5295:5280] * 11301;
    tap_outputs[11695:11680] = value_grid[5311:5296] * 11327;
    tap_outputs[5295:5280] = value_grid[5327:5312] * 11378;
    tap_outputs[5311:5296] = value_grid[5343:5328] * 11430;
    tap_outputs[11743:11728] = value_grid[5359:5344] * 11461;
    tap_outputs[5343:5328] = value_grid[5375:5360] * 11460;
    tap_outputs[11775:11760] = value_grid[5391:5376] * 11429;
    tap_outputs[11791:11776] = value_grid[5407:5392] * 11385;
    tap_outputs[11807:11792] = value_grid[5423:5408] * 11347;
    tap_outputs[5407:5392] = value_grid[5439:5424] * 11330;
    tap_outputs[11839:11824] = value_grid[5455:5440] * 11341;
    tap_outputs[11855:11840] = value_grid[5471:5456] * 11371;
    tap_outputs[11871:11856] = value_grid[5487:5472] * 11407;
    tap_outputs[11887:11872] = value_grid[5503:5488] * 11433;
    tap_outputs[5487:5472] = value_grid[5519:5504] * 11438;
    tap_outputs[11919:11904] = value_grid[5535:5520] * 11423;
    tap_outputs[5519:5504] = value_grid[5551:5536] * 11396;
    tap_outputs[11951:11936] = value_grid[5567:5552] * 11369;
    tap_outputs[11967:11952] = value_grid[5583:5568] * 11353;
    tap_outputs[11983:11968] = value_grid[5599:5584] * 11355;
    tap_outputs[11999:11984] = value_grid[5615:5600] * 11371;
    tap_outputs[5599:5584] = value_grid[5631:5616] * 11394;
    tap_outputs[12031:12016] = value_grid[5647:5632] * 11413;
    tap_outputs[12047:12032] = value_grid[5663:5648] * 11421;
    tap_outputs[12063:12048] = value_grid[5679:5664] * 11415;
    tap_outputs[12079:12064] = value_grid[5695:5680] * 11399;
    tap_outputs[12095:12080] = value_grid[5711:5696] * 11381;
    tap_outputs[12111:12096] = value_grid[5727:5712] * 11369;
    tap_outputs[12127:12112] = value_grid[5743:5728] * 11367;
    tap_outputs[12143:12128] = value_grid[5759:5744] * 11375;
    tap_outputs[5743:5728] = value_grid[5775:5760] * 11388;
    tap_outputs[12175:12160] = value_grid[5791:5776] * 11401;
    tap_outputs[5775:5760] = value_grid[5807:5792] * 11408;
    tap_outputs[12207:12192] = value_grid[5823:5808] * 11407;
    tap_outputs[12223:12208] = value_grid[5839:5824] * 11399;
    tap_outputs[5823:5808] = value_grid[5855:5840] * 11388;
    tap_outputs[5839:5824] = value_grid[5871:5856] * 11380;
    tap_outputs[12271:12256] = value_grid[5887:5872] * 11377;
    tap_outputs[5871:5856] = value_grid[5903:5888] * 11380;
    tap_outputs[12303:12288] = value_grid[5919:5904] * 11387;
    tap_outputs[12319:12304] = value_grid[5935:5920] * 11395;
    tap_outputs[5919:5904] = value_grid[5951:5936] * 11400;
    tap_outputs[5935:5920] = value_grid[5967:5952] * 11400;
    tap_outputs[12367:12352] = value_grid[5983:5968] * 11397;
    tap_outputs[12383:12368] = value_grid[5999:5984] * 11391;
    tap_outputs[5983:5968] = value_grid[6015:6000] * 11386;
    tap_outputs[12415:12400] = value_grid[6031:6016] * 11383;
    tap_outputs[6015:6000] = value_grid[6047:6032] * 11384;
    tap_outputs[12447:12432] = value_grid[6063:6048] * 11387;
    tap_outputs[12463:12448] = value_grid[6079:6064] * 11391;
    tap_outputs[12479:12464] = value_grid[6095:6080] * 11395;
    tap_outputs[6079:6064] = value_grid[6111:6096] * 11396;
    tap_outputs[6095:6080] = value_grid[6127:6112] * 11394;
    tap_outputs[6111:6096] = value_grid[6143:6128] * 11392;
    tap_outputs[12543:12528] = value_grid[6159:6144] * 11389;
    tap_outputs[12559:12544] = value_grid[6175:6160] * 11387;
    tap_outputs[12575:12560] = value_grid[6191:6176] * 11387;
    tap_outputs[6175:6160] = value_grid[6207:6192] * 11388;
    tap_outputs[6191:6176] = value_grid[6223:6208] * 11390;
    tap_outputs[6207:6192] = value_grid[6239:6224] * 11392;
    tap_outputs[12639:12624] = value_grid[6255:6240] * 11393;
    tap_outputs[6239:6224] = value_grid[6271:6256] * 11392;
    tap_outputs[12671:12656] = value_grid[6287:6272] * 11391;
    tap_outputs[6271:6256] = value_grid[6303:6288] * 11390;
    tap_outputs[12703:12688] = value_grid[6319:6304] * 11389;
    tap_outputs[12719:12704] = value_grid[6335:6320] * 11389;
    tap_outputs[12735:12720] = value_grid[6351:6336] * 11389;
    tap_outputs[6335:6320] = value_grid[6367:6352] * 11390;
    tap_outputs[12767:12752] = value_grid[6383:6368] * 11391;
    tap_outputs[12783:12768] = value_grid[6399:6384] * 11391;
    tap_outputs[12799:12784] = value_grid[6415:6400] * 11391;
    tap_outputs[6399:6384] = value_grid[6431:6416] * 11392;
    tap_outputs[6415:6400] = value_grid[6447:6432] * 11390;
    tap_outputs[6431:6416] = value_grid[79:64] * 11390;
    tap_outputs[6447:6432] = value_grid[95:80] * 11392;
    tap_outputs[47:32] = value_grid[111:96] * 11391;
    tap_outputs[63:48] = value_grid[127:112] * 11391;
    tap_outputs[79:64] = value_grid[143:128] * 11391;
    tap_outputs[6511:6496] = value_grid[159:144] * 11390;
    tap_outputs[111:96] = value_grid[175:160] * 11389;
    tap_outputs[127:112] = value_grid[191:176] * 11389;
    tap_outputs[143:128] = value_grid[207:192] * 11389;
    tap_outputs[6575:6560] = value_grid[223:208] * 11390;
    tap_outputs[175:160] = value_grid[239:224] * 11391;
    tap_outputs[6607:6592] = value_grid[255:240] * 11392;
    tap_outputs[207:192] = value_grid[271:256] * 11393;
    tap_outputs[6639:6624] = value_grid[287:272] * 11392;
    tap_outputs[6655:6640] = value_grid[303:288] * 11390;
    tap_outputs[6671:6656] = value_grid[319:304] * 11388;
    tap_outputs[271:256] = value_grid[335:320] * 11387;
    tap_outputs[287:272] = value_grid[351:336] * 11387;
    tap_outputs[303:288] = value_grid[367:352] * 11389;
    tap_outputs[6735:6720] = value_grid[383:368] * 11392;
    tap_outputs[6751:6736] = value_grid[399:384] * 11394;
    tap_outputs[6767:6752] = value_grid[415:400] * 11396;
    tap_outputs[367:352] = value_grid[431:416] * 11395;
    tap_outputs[383:368] = value_grid[447:432] * 11391;
    tap_outputs[399:384] = value_grid[463:448] * 11387;
    tap_outputs[6831:6816] = value_grid[479:464] * 11384;
    tap_outputs[431:416] = value_grid[495:480] * 11383;
    tap_outputs[6863:6848] = value_grid[511:496] * 11386;
    tap_outputs[463:448] = value_grid[527:512] * 11391;
    tap_outputs[479:464] = value_grid[543:528] * 11397;
    tap_outputs[6911:6896] = value_grid[559:544] * 11400;
    tap_outputs[6927:6912] = value_grid[575:560] * 11400;
    tap_outputs[527:512] = value_grid[591:576] * 11395;
    tap_outputs[543:528] = value_grid[607:592] * 11387;
    tap_outputs[6975:6960] = value_grid[623:608] * 11380;
    tap_outputs[575:560] = value_grid[639:624] * 11377;
    tap_outputs[7007:6992] = value_grid[655:640] * 11380;
    tap_outputs[7023:7008] = value_grid[671:656] * 11388;
    tap_outputs[623:608] = value_grid[687:672] * 11399;
    tap_outputs[639:624] = value_grid[703:688] * 11407;
    tap_outputs[7071:7056] = value_grid[719:704] * 11408;
    tap_outputs[671:656] = value_grid[735:720] * 11401;
    tap_outputs[7103:7088] = value_grid[751:736] * 11388;
    tap_outputs[703:688] = value_grid[767:752] * 11375;
    tap_outputs[719:704] = value_grid[783:768] * 11367;
    tap_outputs[735:720] = value_grid[799:784] * 11369;
    tap_outputs[751:736] = value_grid[815:800] * 11381;
    tap_outputs[767:752] = value_grid[831:816] * 11399;
    tap_outputs[783:768] = value_grid[847:832] * 11415;
    tap_outputs[799:784] = value_grid[863:848] * 11421;
    tap_outputs[815:800] = value_grid[879:864] * 11413;
    tap_outputs[7247:7232] = value_grid[895:880] * 11394;
    tap_outputs[847:832] = value_grid[911:896] * 11371;
    tap_outputs[863:848] = value_grid[927:912] * 11355;
    tap_outputs[879:864] = value_grid[943:928] * 11353;
    tap_outputs[895:880] = value_grid[959:944] * 11369;
    tap_outputs[7327:7312] = value_grid[975:960] * 11396;
    tap_outputs[927:912] = value_grid[991:976] * 11423;
    tap_outputs[7359:7344] = value_grid[1007:992] * 11438;
    tap_outputs[959:944] = value_grid[1023:1008] * 11433;
    tap_outputs[975:960] = value_grid[1039:1024] * 11407;
    tap_outputs[991:976] = value_grid[1055:1040] * 11371;
    tap_outputs[1007:992] = value_grid[1071:1056] * 11341;
    tap_outputs[7439:7424] = value_grid[1087:1072] * 11330;
    tap_outputs[1039:1024] = value_grid[1103:1088] * 11347;
    tap_outputs[1055:1040] = value_grid[1119:1104] * 11385;
    tap_outputs[1071:1056] = value_grid[1135:1120] * 11429;
    tap_outputs[7503:7488] = value_grid[1151:1136] * 11460;
    tap_outputs[1103:1088] = value_grid[1167:1152] * 11461;
    tap_outputs[7535:7520] = value_grid[1183:1168] * 11430;
    tap_outputs[7551:7536] = value_grid[1199:1184] * 11378;
    tap_outputs[1151:1136] = value_grid[1215:1200] * 11327;
    tap_outputs[1167:1152] = value_grid[1231:1216] * 11301;
    tap_outputs[7599:7584] = value_grid[1247:1232] * 11314;
    tap_outputs[1199:1184] = value_grid[1263:1248] * 11363;
    tap_outputs[1215:1200] = value_grid[1279:1264] * 11429;
    tap_outputs[1231:1216] = value_grid[1295:1280] * 11483;
    tap_outputs[1247:1232] = value_grid[1311:1296] * 11499;
    tap_outputs[1263:1248] = value_grid[1327:1312] * 11467;
    tap_outputs[7695:7680] = value_grid[1343:1328] * 11396;
    tap_outputs[1295:1280] = value_grid[1359:1344] * 11317;
    tap_outputs[7727:7712] = value_grid[1375:1360] * 11266;
    tap_outputs[1327:1312] = value_grid[1391:1376] * 11267;
    tap_outputs[1343:1328] = value_grid[1407:1392] * 11325;
    tap_outputs[1359:1344] = value_grid[1423:1408] * 11417;
    tap_outputs[1375:1360] = value_grid[1439:1424] * 11505;
    tap_outputs[1391:1376] = value_grid[1455:1440] * 11547;
    tap_outputs[1407:1392] = value_grid[1471:1456] * 11521;
    tap_outputs[1423:1408] = value_grid[1487:1472] * 11433;
    tap_outputs[1439:1424] = value_grid[1503:1488] * 11319;
    tap_outputs[1455:1440] = value_grid[1519:1504] * 11229;
    tap_outputs[7887:7872] = value_grid[1535:1520] * 11206;
    tap_outputs[7903:7888] = value_grid[1551:1536] * 11266;
    tap_outputs[1503:1488] = value_grid[1567:1552] * 11387;
    tap_outputs[1519:1504] = value_grid[1583:1568] * 11519;
    tap_outputs[7951:7936] = value_grid[1599:1584] * 11602;
    tap_outputs[7967:7952] = value_grid[1615:1600] * 11594;
    tap_outputs[1567:1552] = value_grid[1631:1616] * 11493;
    tap_outputs[7999:7984] = value_grid[1647:1632] * 11338;
    tap_outputs[8015:8000] = value_grid[1663:1648] * 11196;
    tap_outputs[8031:8016] = value_grid[1679:1664] * 11132;
    tap_outputs[1631:1616] = value_grid[1695:1680] * 11181;
    tap_outputs[8063:8048] = value_grid[1711:1696] * 11330;
    tap_outputs[8079:8064] = value_grid[1727:1712] * 11516;
    tap_outputs[8095:8080] = value_grid[1743:1728] * 11658;
    tap_outputs[8111:8096] = value_grid[1759:1744] * 11688;
    tap_outputs[8127:8112] = value_grid[1775:1760] * 11584;
    tap_outputs[8143:8128] = value_grid[1791:1776] * 11386;
    tap_outputs[8159:8144] = value_grid[1807:1792] * 11176;
    tap_outputs[1759:1744] = value_grid[1823:1808] * 11049;
    tap_outputs[1775:1760] = value_grid[1839:1824] * 11069;
    tap_outputs[1791:1776] = value_grid[1855:1840] * 11237;
    tap_outputs[1807:1792] = value_grid[1871:1856] * 11485;
    tap_outputs[1823:1808] = value_grid[1887:1872] * 11707;
    tap_outputs[1839:1824] = value_grid[1903:1888] * 11799;
    tap_outputs[8271:8256] = value_grid[1919:1904] * 11712;
    tap_outputs[1871:1856] = value_grid[1935:1920] * 11473;
    tap_outputs[8303:8288] = value_grid[1951:1936] * 11180;
    tap_outputs[1903:1888] = value_grid[1967:1952] * 10965;
    tap_outputs[1919:1904] = value_grid[1983:1968] * 10929;
    tap_outputs[8351:8336] = value_grid[1999:1984] * 11100;
    tap_outputs[8367:8352] = value_grid[2015:2000] * 11414;
    tap_outputs[1967:1952] = value_grid[2031:2016] * 11737;
    tap_outputs[8399:8384] = value_grid[2047:2032] * 11924;
    tap_outputs[8415:8400] = value_grid[2063:2048] * 11880;
    tap_outputs[2015:2000] = value_grid[2079:2064] * 11611;
    tap_outputs[2031:2016] = value_grid[2095:2080] * 11225;
    tap_outputs[2047:2032] = value_grid[2111:2096] * 10891;
    tap_outputs[2063:2048] = value_grid[2127:2112] * 10761;
    tap_outputs[8495:8480] = value_grid[2143:2128] * 10910;
    tap_outputs[2095:2080] = value_grid[2159:2144] * 11285;
    tap_outputs[2111:2096] = value_grid[2175:2160] * 11731;
    tap_outputs[2127:2112] = value_grid[2191:2176] * 12051;
    tap_outputs[8559:8544] = value_grid[2207:2192] * 12090;
    tap_outputs[2159:2144] = value_grid[2223:2208] * 11815;
    tap_outputs[8591:8576] = value_grid[2239:2224] * 11330;
    tap_outputs[8607:8592] = value_grid[2255:2240] * 10842;
    tap_outputs[2207:2192] = value_grid[2271:2256] * 10573;
    tap_outputs[8639:8624] = value_grid[2287:2272] * 10658;
    tap_outputs[8655:8640] = value_grid[2303:2288] * 11080;
    tap_outputs[2255:2240] = value_grid[2319:2304] * 11669;
    tap_outputs[8687:8672] = value_grid[2335:2320] * 12168;
    tap_outputs[2287:2272] = value_grid[2351:2336] * 12345;
    tap_outputs[2303:2288] = value_grid[2367:2352] * 12101;
    tap_outputs[2319:2304] = value_grid[2383:2368] * 11519;
    tap_outputs[8751:8736] = value_grid[2399:2384] * 10842;
    tap_outputs[8767:8752] = value_grid[2415:2400] * 10372;
    tap_outputs[8783:8768] = value_grid[2431:2416] * 10334;
    tap_outputs[2383:2368] = value_grid[2447:2432] * 10773;
    tap_outputs[8815:8800] = value_grid[2463:2448] * 11520;
    tap_outputs[2415:2400] = value_grid[2479:2464] * 12255;
    tap_outputs[2431:2416] = value_grid[2495:2480] * 12645;
    tap_outputs[8863:8848] = value_grid[2511:2496] * 12490;
    tap_outputs[8879:8864] = value_grid[2527:2512] * 11826;
    tap_outputs[2479:2464] = value_grid[2543:2528] * 10921;
    tap_outputs[8911:8896] = value_grid[2559:2544] * 10170;
    tap_outputs[2511:2496] = value_grid[2575:2560] * 9923;
    tap_outputs[2527:2512] = value_grid[2591:2576] * 10327;
    tap_outputs[2543:2528] = value_grid[2607:2592] * 11241;
    tap_outputs[2559:2544] = value_grid[2623:2608] * 12285;
    tap_outputs[2575:2560] = value_grid[2639:2624] * 12995;
    tap_outputs[2591:2576] = value_grid[2655:2640] * 13023;
    tap_outputs[2607:2592] = value_grid[2671:2656] * 12311;
    tap_outputs[9039:9024] = value_grid[2687:2672] * 11128;
    tap_outputs[2639:2624] = value_grid[2703:2688] * 9979;
    tap_outputs[9071:9056] = value_grid[2719:2704] * 9388;
    tap_outputs[2671:2656] = value_grid[2735:2720] * 9667;
    tap_outputs[9103:9088] = value_grid[2751:2736] * 10754;
    tap_outputs[9119:9104] = value_grid[2767:2752] * 12216;
    tap_outputs[9135:9120] = value_grid[2783:2768] * 13416;
    tap_outputs[2735:2720] = value_grid[2799:2784] * 13787;
    tap_outputs[2751:2736] = value_grid[2815:2800] * 13091;
    tap_outputs[2767:2752] = value_grid[2831:2816] * 11557;
    tap_outputs[9199:9184] = value_grid[2847:2832] * 9812;
    tap_outputs[2799:2784] = value_grid[2863:2848] * 8637;
    tap_outputs[2815:2800] = value_grid[2879:2864] * 8619;
    tap_outputs[2831:2816] = value_grid[2895:2880] * 9877;
    tap_outputs[9263:9248] = value_grid[2911:2896] * 11956;
    tap_outputs[2863:2848] = value_grid[2927:2912] * 13985;
    tap_outputs[9295:9280] = value_grid[2943:2928] * 15028;
    tap_outputs[9311:9296] = value_grid[2959:2944] * 14498;
    tap_outputs[2911:2896] = value_grid[2975:2960] * 12463;
    tap_outputs[2927:2912] = value_grid[2991:2976] * 9683;
    tap_outputs[9359:9344] = value_grid[3007:2992] * 7350;
    tap_outputs[9375:9360] = value_grid[3023:3008] * 6602;
    tap_outputs[2975:2960] = value_grid[3039:3024] * 8001;
    tap_outputs[2991:2976] = value_grid[3055:3040] * 11213;
    tap_outputs[9423:9408] = value_grid[3071:3056] * 15026;
    tap_outputs[9439:9424] = value_grid[3087:3072] * 17762;
    tap_outputs[3039:3024] = value_grid[3103:3088] * 17947;
    tap_outputs[9471:9456] = value_grid[3119:3104] * 14992;
    tap_outputs[3071:3056] = value_grid[3135:3120] * 9601;
    tap_outputs[3087:3072] = value_grid[3151:3136] * 3723;
    tap_outputs[9519:9504] = value_grid[3167:3152] * 0;
    tap_outputs[9535:9520] = value_grid[3183:3168] * 874;
    tap_outputs[3135:3120] = value_grid[3199:3184] * 7657;
    tap_outputs[3151:3136] = value_grid[3215:3200] * 19907;
    tap_outputs[9583:9568] = value_grid[3231:3216] * 35362;
    tap_outputs[3183:3168] = value_grid[3247:3232] * 50489;
    tap_outputs[3199:3184] = value_grid[3263:3248] * 61505;
    tap_outputs[3215:3200] = value_grid[3279:3264] * 65535;
    tap_outputs[3231:3216] = value_grid[3295:3280] * 61505;
    tap_outputs[3247:3232] = value_grid[3311:3296] * 50489;
    tap_outputs[9679:9664] = value_grid[3327:3312] * 35362;
    tap_outputs[3279:3264] = value_grid[3343:3328] * 19907;
    tap_outputs[3295:3280] = value_grid[3359:3344] * 7657;
    tap_outputs[9727:9712] = value_grid[3375:3360] * 874;
    tap_outputs[9743:9728] = value_grid[3391:3376] * 0;
    tap_outputs[3343:3328] = value_grid[3407:3392] * 3723;
    tap_outputs[3359:3344] = value_grid[3423:3408] * 9601;
    tap_outputs[9791:9776] = value_grid[3439:3424] * 14992;
    tap_outputs[3391:3376] = value_grid[3455:3440] * 17947;
    tap_outputs[9823:9808] = value_grid[3471:3456] * 17762;
    tap_outputs[9839:9824] = value_grid[3487:3472] * 15026;
    tap_outputs[3439:3424] = value_grid[3503:3488] * 11213;
    tap_outputs[3455:3440] = value_grid[3519:3504] * 8001;
    tap_outputs[9887:9872] = value_grid[3535:3520] * 6602;
    tap_outputs[9903:9888] = value_grid[3551:3536] * 7350;
    tap_outputs[3503:3488] = value_grid[3567:3552] * 9683;
    tap_outputs[3519:3504] = value_grid[3583:3568] * 12463;
    tap_outputs[9951:9936] = value_grid[3599:3584] * 14498;
    tap_outputs[9967:9952] = value_grid[3615:3600] * 15028;
    tap_outputs[3567:3552] = value_grid[3631:3616] * 13985;
    tap_outputs[9999:9984] = value_grid[3647:3632] * 11956;
    tap_outputs[3599:3584] = value_grid[3663:3648] * 9877;
    tap_outputs[3615:3600] = value_grid[3679:3664] * 8619;
    tap_outputs[3631:3616] = value_grid[3695:3680] * 8637;
    tap_outputs[10063:10048] = value_grid[3711:3696] * 9812;
    tap_outputs[3663:3648] = value_grid[3727:3712] * 11557;
    tap_outputs[3679:3664] = value_grid[3743:3728] * 13091;
    tap_outputs[3695:3680] = value_grid[3759:3744] * 13787;
    tap_outputs[10127:10112] = value_grid[3775:3760] * 13416;
    tap_outputs[10143:10128] = value_grid[3791:3776] * 12216;
    tap_outputs[10159:10144] = value_grid[3807:3792] * 10754;
    tap_outputs[3759:3744] = value_grid[3823:3808] * 9667;
    tap_outputs[10191:10176] = value_grid[3839:3824] * 9388;
    tap_outputs[3791:3776] = value_grid[3855:3840] * 9979;
    tap_outputs[10223:10208] = value_grid[3871:3856] * 11128;
    tap_outputs[3823:3808] = value_grid[3887:3872] * 12311;
    tap_outputs[3839:3824] = value_grid[3903:3888] * 13023;
    tap_outputs[3855:3840] = value_grid[3919:3904] * 12995;
    tap_outputs[3871:3856] = value_grid[3935:3920] * 12285;
    tap_outputs[3887:3872] = value_grid[3951:3936] * 11241;
    tap_outputs[3903:3888] = value_grid[3967:3952] * 10327;
    tap_outputs[3919:3904] = value_grid[3983:3968] * 9923;
    tap_outputs[10351:10336] = value_grid[3999:3984] * 10170;
    tap_outputs[3951:3936] = value_grid[4015:4000] * 10921;
    tap_outputs[10383:10368] = value_grid[4031:4016] * 11826;
    tap_outputs[10399:10384] = value_grid[4047:4032] * 12490;
    tap_outputs[3999:3984] = value_grid[4063:4048] * 12645;
    tap_outputs[4015:4000] = value_grid[4079:4064] * 12255;
    tap_outputs[10447:10432] = value_grid[4095:4080] * 11520;
    tap_outputs[4047:4032] = value_grid[4111:4096] * 10773;
    tap_outputs[10479:10464] = value_grid[4127:4112] * 10334;
    tap_outputs[10495:10480] = value_grid[4143:4128] * 10372;
    tap_outputs[10511:10496] = value_grid[4159:4144] * 10842;
    tap_outputs[4111:4096] = value_grid[4175:4160] * 11519;
    tap_outputs[4127:4112] = value_grid[4191:4176] * 12101;
    tap_outputs[4143:4128] = value_grid[4207:4192] * 12345;
    tap_outputs[10575:10560] = value_grid[4223:4208] * 12168;
    tap_outputs[4175:4160] = value_grid[4239:4224] * 11669;
    tap_outputs[10607:10592] = value_grid[4255:4240] * 11080;
    tap_outputs[10623:10608] = value_grid[4271:4256] * 10658;
    tap_outputs[4223:4208] = value_grid[4287:4272] * 10573;
    tap_outputs[10655:10640] = value_grid[4303:4288] * 10842;
    tap_outputs[10671:10656] = value_grid[4319:4304] * 11330;
    tap_outputs[4271:4256] = value_grid[4335:4320] * 11815;
    tap_outputs[10703:10688] = value_grid[4351:4336] * 12090;
    tap_outputs[4303:4288] = value_grid[4367:4352] * 12051;
    tap_outputs[4319:4304] = value_grid[4383:4368] * 11731;
    tap_outputs[4335:4320] = value_grid[4399:4384] * 11285;
    tap_outputs[10767:10752] = value_grid[4415:4400] * 10910;
    tap_outputs[4367:4352] = value_grid[4431:4416] * 10761;
    tap_outputs[4383:4368] = value_grid[4447:4432] * 10891;
    tap_outputs[4399:4384] = value_grid[4463:4448] * 11225;
    tap_outputs[4415:4400] = value_grid[4479:4464] * 11611;
    tap_outputs[10847:10832] = value_grid[4495:4480] * 11880;
    tap_outputs[10863:10848] = value_grid[4511:4496] * 11924;
    tap_outputs[4463:4448] = value_grid[4527:4512] * 11737;
    tap_outputs[10895:10880] = value_grid[4543:4528] * 11414;
    tap_outputs[10911:10896] = value_grid[4559:4544] * 11100;
    tap_outputs[4511:4496] = value_grid[4575:4560] * 10929;
    tap_outputs[4527:4512] = value_grid[4591:4576] * 10965;
    tap_outputs[10959:10944] = value_grid[4607:4592] * 11180;
    tap_outputs[4559:4544] = value_grid[4623:4608] * 11473;
    tap_outputs[10991:10976] = value_grid[4639:4624] * 11712;
    tap_outputs[4591:4576] = value_grid[4655:4640] * 11799;
    tap_outputs[4607:4592] = value_grid[4671:4656] * 11707;
    tap_outputs[4623:4608] = value_grid[4687:4672] * 11485;
    tap_outputs[4639:4624] = value_grid[4703:4688] * 11237;
    tap_outputs[4655:4640] = value_grid[4719:4704] * 11069;
    tap_outputs[4671:4656] = value_grid[4735:4720] * 11049;
    tap_outputs[11103:11088] = value_grid[4751:4736] * 11176;
    tap_outputs[11119:11104] = value_grid[4767:4752] * 11386;
    tap_outputs[11135:11120] = value_grid[4783:4768] * 11584;
    tap_outputs[11151:11136] = value_grid[4799:4784] * 11688;
    tap_outputs[11167:11152] = value_grid[4815:4800] * 11658;
    tap_outputs[11183:11168] = value_grid[4831:4816] * 11516;
    tap_outputs[11199:11184] = value_grid[4847:4832] * 11330;
    tap_outputs[4799:4784] = value_grid[4863:4848] * 11181;
    tap_outputs[11231:11216] = value_grid[4879:4864] * 11132;
    tap_outputs[11247:11232] = value_grid[4895:4880] * 11196;
    tap_outputs[11263:11248] = value_grid[4911:4896] * 11338;
    tap_outputs[4863:4848] = value_grid[4927:4912] * 11493;
    tap_outputs[11295:11280] = value_grid[4943:4928] * 11594;
    tap_outputs[11311:11296] = value_grid[4959:4944] * 11602;
    tap_outputs[4911:4896] = value_grid[4975:4960] * 11519;
    tap_outputs[4927:4912] = value_grid[4991:4976] * 11387;
    tap_outputs[11359:11344] = value_grid[5007:4992] * 11266;
    tap_outputs[11375:11360] = value_grid[5023:5008] * 11206;
    tap_outputs[4975:4960] = value_grid[5039:5024] * 11229;
    tap_outputs[4991:4976] = value_grid[5055:5040] * 11319;
    tap_outputs[5007:4992] = value_grid[5071:5056] * 11433;
    tap_outputs[5023:5008] = value_grid[5087:5072] * 11521;
    tap_outputs[5039:5024] = value_grid[5103:5088] * 11547;
    tap_outputs[5055:5040] = value_grid[5119:5104] * 11505;
    tap_outputs[5071:5056] = value_grid[5135:5120] * 11417;
    tap_outputs[5087:5072] = value_grid[5151:5136] * 11325;
    tap_outputs[5103:5088] = value_grid[5167:5152] * 11267;
    tap_outputs[11535:11520] = value_grid[5183:5168] * 11266;
    tap_outputs[5135:5120] = value_grid[5199:5184] * 11317;
    tap_outputs[11567:11552] = value_grid[5215:5200] * 11396;
    tap_outputs[5167:5152] = value_grid[5231:5216] * 11467;
    tap_outputs[5183:5168] = value_grid[5247:5232] * 11499;
    tap_outputs[5199:5184] = value_grid[5263:5248] * 11483;
    tap_outputs[5215:5200] = value_grid[5279:5264] * 11429;
    tap_outputs[5231:5216] = value_grid[5295:5280] * 11363;
    tap_outputs[11663:11648] = value_grid[5311:5296] * 11314;
    tap_outputs[5263:5248] = value_grid[5327:5312] * 11301;
    tap_outputs[5279:5264] = value_grid[5343:5328] * 11327;
    tap_outputs[11711:11696] = value_grid[5359:5344] * 11378;
    tap_outputs[11727:11712] = value_grid[5375:5360] * 11430;
    tap_outputs[5327:5312] = value_grid[5391:5376] * 11461;
    tap_outputs[11759:11744] = value_grid[5407:5392] * 11460;
    tap_outputs[5359:5344] = value_grid[5423:5408] * 11429;
    tap_outputs[5375:5360] = value_grid[5439:5424] * 11385;
    tap_outputs[5391:5376] = value_grid[5455:5440] * 11347;
    tap_outputs[11823:11808] = value_grid[5471:5456] * 11330;
    tap_outputs[5423:5408] = value_grid[5487:5472] * 11341;
    tap_outputs[5439:5424] = value_grid[5503:5488] * 11371;
    tap_outputs[5455:5440] = value_grid[5519:5504] * 11407;
    tap_outputs[5471:5456] = value_grid[5535:5520] * 11433;
    tap_outputs[11903:11888] = value_grid[5551:5536] * 11438;
    tap_outputs[5503:5488] = value_grid[5567:5552] * 11423;
    tap_outputs[11935:11920] = value_grid[5583:5568] * 11396;
    tap_outputs[5535:5520] = value_grid[5599:5584] * 11369;
    tap_outputs[5551:5536] = value_grid[5615:5600] * 11353;
    tap_outputs[5567:5552] = value_grid[5631:5616] * 11355;
    tap_outputs[5583:5568] = value_grid[5647:5632] * 11371;
    tap_outputs[12015:12000] = value_grid[5663:5648] * 11394;
    tap_outputs[5615:5600] = value_grid[5679:5664] * 11413;
    tap_outputs[5631:5616] = value_grid[5695:5680] * 11421;
    tap_outputs[5647:5632] = value_grid[5711:5696] * 11415;
    tap_outputs[5663:5648] = value_grid[5727:5712] * 11399;
    tap_outputs[5679:5664] = value_grid[5743:5728] * 11381;
    tap_outputs[5695:5680] = value_grid[5759:5744] * 11369;
    tap_outputs[5711:5696] = value_grid[5775:5760] * 11367;
    tap_outputs[5727:5712] = value_grid[5791:5776] * 11375;
    tap_outputs[12159:12144] = value_grid[5807:5792] * 11388;
    tap_outputs[5759:5744] = value_grid[5823:5808] * 11401;
    tap_outputs[12191:12176] = value_grid[5839:5824] * 11408;
    tap_outputs[5791:5776] = value_grid[5855:5840] * 11407;
    tap_outputs[5807:5792] = value_grid[5871:5856] * 11399;
    tap_outputs[12239:12224] = value_grid[5887:5872] * 11388;
    tap_outputs[12255:12240] = value_grid[5903:5888] * 11380;
    tap_outputs[5855:5840] = value_grid[5919:5904] * 11377;
    tap_outputs[12287:12272] = value_grid[5935:5920] * 11380;
    tap_outputs[5887:5872] = value_grid[5951:5936] * 11387;
    tap_outputs[5903:5888] = value_grid[5967:5952] * 11395;
    tap_outputs[12335:12320] = value_grid[5983:5968] * 11400;
    tap_outputs[12351:12336] = value_grid[5999:5984] * 11400;
    tap_outputs[5951:5936] = value_grid[6015:6000] * 11397;
    tap_outputs[5967:5952] = value_grid[6031:6016] * 11391;
    tap_outputs[12399:12384] = value_grid[6047:6032] * 11386;
    tap_outputs[5999:5984] = value_grid[6063:6048] * 11383;
    tap_outputs[12431:12416] = value_grid[6079:6064] * 11384;
    tap_outputs[6031:6016] = value_grid[6095:6080] * 11387;
    tap_outputs[6047:6032] = value_grid[6111:6096] * 11391;
    tap_outputs[6063:6048] = value_grid[6127:6112] * 11395;
    tap_outputs[12495:12480] = value_grid[6143:6128] * 11396;
    tap_outputs[12511:12496] = value_grid[6159:6144] * 11394;
    tap_outputs[12527:12512] = value_grid[6175:6160] * 11392;
    tap_outputs[6127:6112] = value_grid[6191:6176] * 11389;
    tap_outputs[6143:6128] = value_grid[6207:6192] * 11387;
    tap_outputs[6159:6144] = value_grid[6223:6208] * 11387;
    tap_outputs[12591:12576] = value_grid[6239:6224] * 11388;
    tap_outputs[12607:12592] = value_grid[6255:6240] * 11390;
    tap_outputs[12623:12608] = value_grid[6271:6256] * 11392;
    tap_outputs[6223:6208] = value_grid[6287:6272] * 11393;
    tap_outputs[12655:12640] = value_grid[6303:6288] * 11392;
    tap_outputs[6255:6240] = value_grid[6319:6304] * 11391;
    tap_outputs[12687:12672] = value_grid[6335:6320] * 11390;
    tap_outputs[6287:6272] = value_grid[6351:6336] * 11389;
    tap_outputs[6303:6288] = value_grid[6367:6352] * 11389;
    tap_outputs[6319:6304] = value_grid[6383:6368] * 11389;
    tap_outputs[12751:12736] = value_grid[6399:6384] * 11390;
    tap_outputs[6351:6336] = value_grid[6415:6400] * 11391;
    tap_outputs[6367:6352] = value_grid[6431:6416] * 11391;
    tap_outputs[6383:6368] = value_grid[6447:6432] * 11391;
    tap_outputs[12815:12800] = value_grid[6463:6448] * 11392;
    tap_outputs[12831:12816] = value_grid[6479:6464] * 11390;
    adder_tree_tier_0_p0_in = tap_outputs[6415:0];
    adder_tree_tier_1_p0_in[15:0] = adder_tree_tier_0_p0_in[15:0] + adder_tree_tier_0_p0_in[31:16];
    adder_tree_tier_1_p0_in[31:16] = adder_tree_tier_0_p0_in[47:32] + adder_tree_tier_0_p0_in[63:48];
    adder_tree_tier_1_p0_in[47:32] = adder_tree_tier_0_p0_in[79:64] + adder_tree_tier_0_p0_in[95:80];
    adder_tree_tier_1_p0_in[63:48] = adder_tree_tier_0_p0_in[111:96] + adder_tree_tier_0_p0_in[127:112];
    adder_tree_tier_1_p0_in[79:64] = adder_tree_tier_0_p0_in[143:128] + adder_tree_tier_0_p0_in[159:144];
    adder_tree_tier_1_p0_in[95:80] = adder_tree_tier_0_p0_in[175:160] + adder_tree_tier_0_p0_in[191:176];
    adder_tree_tier_1_p0_in[111:96] = adder_tree_tier_0_p0_in[207:192] + adder_tree_tier_0_p0_in[223:208];
    adder_tree_tier_1_p0_in[127:112] = adder_tree_tier_0_p0_in[239:224] + adder_tree_tier_0_p0_in[255:240];
    adder_tree_tier_1_p0_in[143:128] = adder_tree_tier_0_p0_in[271:256] + adder_tree_tier_0_p0_in[287:272];
    adder_tree_tier_1_p0_in[159:144] = adder_tree_tier_0_p0_in[303:288] + adder_tree_tier_0_p0_in[319:304];
    adder_tree_tier_1_p0_in[175:160] = adder_tree_tier_0_p0_in[335:320] + adder_tree_tier_0_p0_in[351:336];
    adder_tree_tier_1_p0_in[191:176] = adder_tree_tier_0_p0_in[367:352] + adder_tree_tier_0_p0_in[383:368];
    adder_tree_tier_1_p0_in[207:192] = adder_tree_tier_0_p0_in[399:384] + adder_tree_tier_0_p0_in[415:400];
    adder_tree_tier_1_p0_in[223:208] = adder_tree_tier_0_p0_in[431:416] + adder_tree_tier_0_p0_in[447:432];
    adder_tree_tier_1_p0_in[239:224] = adder_tree_tier_0_p0_in[463:448] + adder_tree_tier_0_p0_in[479:464];
    adder_tree_tier_1_p0_in[255:240] = adder_tree_tier_0_p0_in[495:480] + adder_tree_tier_0_p0_in[511:496];
    adder_tree_tier_1_p0_in[271:256] = adder_tree_tier_0_p0_in[527:512] + adder_tree_tier_0_p0_in[543:528];
    adder_tree_tier_1_p0_in[287:272] = adder_tree_tier_0_p0_in[559:544] + adder_tree_tier_0_p0_in[575:560];
    adder_tree_tier_1_p0_in[303:288] = adder_tree_tier_0_p0_in[591:576] + adder_tree_tier_0_p0_in[607:592];
    adder_tree_tier_1_p0_in[319:304] = adder_tree_tier_0_p0_in[623:608] + adder_tree_tier_0_p0_in[639:624];
    adder_tree_tier_1_p0_in[335:320] = adder_tree_tier_0_p0_in[655:640] + adder_tree_tier_0_p0_in[671:656];
    adder_tree_tier_1_p0_in[351:336] = adder_tree_tier_0_p0_in[687:672] + adder_tree_tier_0_p0_in[703:688];
    adder_tree_tier_1_p0_in[367:352] = adder_tree_tier_0_p0_in[719:704] + adder_tree_tier_0_p0_in[735:720];
    adder_tree_tier_1_p0_in[383:368] = adder_tree_tier_0_p0_in[751:736] + adder_tree_tier_0_p0_in[767:752];
    adder_tree_tier_1_p0_in[399:384] = adder_tree_tier_0_p0_in[783:768] + adder_tree_tier_0_p0_in[799:784];
    adder_tree_tier_1_p0_in[415:400] = adder_tree_tier_0_p0_in[815:800] + adder_tree_tier_0_p0_in[831:816];
    adder_tree_tier_1_p0_in[431:416] = adder_tree_tier_0_p0_in[847:832] + adder_tree_tier_0_p0_in[863:848];
    adder_tree_tier_1_p0_in[447:432] = adder_tree_tier_0_p0_in[879:864] + adder_tree_tier_0_p0_in[895:880];
    adder_tree_tier_1_p0_in[463:448] = adder_tree_tier_0_p0_in[911:896] + adder_tree_tier_0_p0_in[927:912];
    adder_tree_tier_1_p0_in[479:464] = adder_tree_tier_0_p0_in[943:928] + adder_tree_tier_0_p0_in[959:944];
    adder_tree_tier_1_p0_in[495:480] = adder_tree_tier_0_p0_in[975:960] + adder_tree_tier_0_p0_in[991:976];
    adder_tree_tier_1_p0_in[511:496] = adder_tree_tier_0_p0_in[1007:992] + adder_tree_tier_0_p0_in[1023:1008];
    adder_tree_tier_1_p0_in[527:512] = adder_tree_tier_0_p0_in[1039:1024] + adder_tree_tier_0_p0_in[1055:1040];
    adder_tree_tier_1_p0_in[543:528] = adder_tree_tier_0_p0_in[1071:1056] + adder_tree_tier_0_p0_in[1087:1072];
    adder_tree_tier_1_p0_in[559:544] = adder_tree_tier_0_p0_in[1103:1088] + adder_tree_tier_0_p0_in[1119:1104];
    adder_tree_tier_1_p0_in[575:560] = adder_tree_tier_0_p0_in[1135:1120] + adder_tree_tier_0_p0_in[1151:1136];
    adder_tree_tier_1_p0_in[591:576] = adder_tree_tier_0_p0_in[1167:1152] + adder_tree_tier_0_p0_in[1183:1168];
    adder_tree_tier_1_p0_in[607:592] = adder_tree_tier_0_p0_in[1199:1184] + adder_tree_tier_0_p0_in[1215:1200];
    adder_tree_tier_1_p0_in[623:608] = adder_tree_tier_0_p0_in[1231:1216] + adder_tree_tier_0_p0_in[1247:1232];
    adder_tree_tier_1_p0_in[639:624] = adder_tree_tier_0_p0_in[1263:1248] + adder_tree_tier_0_p0_in[1279:1264];
    adder_tree_tier_1_p0_in[655:640] = adder_tree_tier_0_p0_in[1295:1280] + adder_tree_tier_0_p0_in[1311:1296];
    adder_tree_tier_1_p0_in[671:656] = adder_tree_tier_0_p0_in[1327:1312] + adder_tree_tier_0_p0_in[1343:1328];
    adder_tree_tier_1_p0_in[687:672] = adder_tree_tier_0_p0_in[1359:1344] + adder_tree_tier_0_p0_in[1375:1360];
    adder_tree_tier_1_p0_in[703:688] = adder_tree_tier_0_p0_in[1391:1376] + adder_tree_tier_0_p0_in[1407:1392];
    adder_tree_tier_1_p0_in[719:704] = adder_tree_tier_0_p0_in[1423:1408] + adder_tree_tier_0_p0_in[1439:1424];
    adder_tree_tier_1_p0_in[735:720] = adder_tree_tier_0_p0_in[1455:1440] + adder_tree_tier_0_p0_in[1471:1456];
    adder_tree_tier_1_p0_in[751:736] = adder_tree_tier_0_p0_in[1487:1472] + adder_tree_tier_0_p0_in[1503:1488];
    adder_tree_tier_1_p0_in[767:752] = adder_tree_tier_0_p0_in[1519:1504] + adder_tree_tier_0_p0_in[1535:1520];
    adder_tree_tier_1_p0_in[783:768] = adder_tree_tier_0_p0_in[1551:1536] + adder_tree_tier_0_p0_in[1567:1552];
    adder_tree_tier_1_p0_in[799:784] = adder_tree_tier_0_p0_in[1583:1568] + adder_tree_tier_0_p0_in[1599:1584];
    adder_tree_tier_1_p0_in[815:800] = adder_tree_tier_0_p0_in[1615:1600] + adder_tree_tier_0_p0_in[1631:1616];
    adder_tree_tier_1_p0_in[831:816] = adder_tree_tier_0_p0_in[1647:1632] + adder_tree_tier_0_p0_in[1663:1648];
    adder_tree_tier_1_p0_in[847:832] = adder_tree_tier_0_p0_in[1679:1664] + adder_tree_tier_0_p0_in[1695:1680];
    adder_tree_tier_1_p0_in[863:848] = adder_tree_tier_0_p0_in[1711:1696] + adder_tree_tier_0_p0_in[1727:1712];
    adder_tree_tier_1_p0_in[879:864] = adder_tree_tier_0_p0_in[1743:1728] + adder_tree_tier_0_p0_in[1759:1744];
    adder_tree_tier_1_p0_in[895:880] = adder_tree_tier_0_p0_in[1775:1760] + adder_tree_tier_0_p0_in[1791:1776];
    adder_tree_tier_1_p0_in[911:896] = adder_tree_tier_0_p0_in[1807:1792] + adder_tree_tier_0_p0_in[1823:1808];
    adder_tree_tier_1_p0_in[927:912] = adder_tree_tier_0_p0_in[1839:1824] + adder_tree_tier_0_p0_in[1855:1840];
    adder_tree_tier_1_p0_in[943:928] = adder_tree_tier_0_p0_in[1871:1856] + adder_tree_tier_0_p0_in[1887:1872];
    adder_tree_tier_1_p0_in[959:944] = adder_tree_tier_0_p0_in[1903:1888] + adder_tree_tier_0_p0_in[1919:1904];
    adder_tree_tier_1_p0_in[975:960] = adder_tree_tier_0_p0_in[1935:1920] + adder_tree_tier_0_p0_in[1951:1936];
    adder_tree_tier_1_p0_in[991:976] = adder_tree_tier_0_p0_in[1967:1952] + adder_tree_tier_0_p0_in[1983:1968];
    adder_tree_tier_1_p0_in[1007:992] = adder_tree_tier_0_p0_in[1999:1984] + adder_tree_tier_0_p0_in[2015:2000];
    adder_tree_tier_1_p0_in[1023:1008] = adder_tree_tier_0_p0_in[2031:2016] + adder_tree_tier_0_p0_in[2047:2032];
    adder_tree_tier_1_p0_in[1039:1024] = adder_tree_tier_0_p0_in[2063:2048] + adder_tree_tier_0_p0_in[2079:2064];
    adder_tree_tier_1_p0_in[1055:1040] = adder_tree_tier_0_p0_in[2095:2080] + adder_tree_tier_0_p0_in[2111:2096];
    adder_tree_tier_1_p0_in[1071:1056] = adder_tree_tier_0_p0_in[2127:2112] + adder_tree_tier_0_p0_in[2143:2128];
    adder_tree_tier_1_p0_in[1087:1072] = adder_tree_tier_0_p0_in[2159:2144] + adder_tree_tier_0_p0_in[2175:2160];
    adder_tree_tier_1_p0_in[1103:1088] = adder_tree_tier_0_p0_in[2191:2176] + adder_tree_tier_0_p0_in[2207:2192];
    adder_tree_tier_1_p0_in[1119:1104] = adder_tree_tier_0_p0_in[2223:2208] + adder_tree_tier_0_p0_in[2239:2224];
    adder_tree_tier_1_p0_in[1135:1120] = adder_tree_tier_0_p0_in[2255:2240] + adder_tree_tier_0_p0_in[2271:2256];
    adder_tree_tier_1_p0_in[1151:1136] = adder_tree_tier_0_p0_in[2287:2272] + adder_tree_tier_0_p0_in[2303:2288];
    adder_tree_tier_1_p0_in[1167:1152] = adder_tree_tier_0_p0_in[2319:2304] + adder_tree_tier_0_p0_in[2335:2320];
    adder_tree_tier_1_p0_in[1183:1168] = adder_tree_tier_0_p0_in[2351:2336] + adder_tree_tier_0_p0_in[2367:2352];
    adder_tree_tier_1_p0_in[1199:1184] = adder_tree_tier_0_p0_in[2383:2368] + adder_tree_tier_0_p0_in[2399:2384];
    adder_tree_tier_1_p0_in[1215:1200] = adder_tree_tier_0_p0_in[2415:2400] + adder_tree_tier_0_p0_in[2431:2416];
    adder_tree_tier_1_p0_in[1231:1216] = adder_tree_tier_0_p0_in[2447:2432] + adder_tree_tier_0_p0_in[2463:2448];
    adder_tree_tier_1_p0_in[1247:1232] = adder_tree_tier_0_p0_in[2479:2464] + adder_tree_tier_0_p0_in[2495:2480];
    adder_tree_tier_1_p0_in[1263:1248] = adder_tree_tier_0_p0_in[2511:2496] + adder_tree_tier_0_p0_in[2527:2512];
    adder_tree_tier_1_p0_in[1279:1264] = adder_tree_tier_0_p0_in[2543:2528] + adder_tree_tier_0_p0_in[2559:2544];
    adder_tree_tier_1_p0_in[1295:1280] = adder_tree_tier_0_p0_in[2575:2560] + adder_tree_tier_0_p0_in[2591:2576];
    adder_tree_tier_1_p0_in[1311:1296] = adder_tree_tier_0_p0_in[2607:2592] + adder_tree_tier_0_p0_in[2623:2608];
    adder_tree_tier_1_p0_in[1327:1312] = adder_tree_tier_0_p0_in[2639:2624] + adder_tree_tier_0_p0_in[2655:2640];
    adder_tree_tier_1_p0_in[1343:1328] = adder_tree_tier_0_p0_in[2671:2656] + adder_tree_tier_0_p0_in[2687:2672];
    adder_tree_tier_1_p0_in[1359:1344] = adder_tree_tier_0_p0_in[2703:2688] + adder_tree_tier_0_p0_in[2719:2704];
    adder_tree_tier_1_p0_in[1375:1360] = adder_tree_tier_0_p0_in[2735:2720] + adder_tree_tier_0_p0_in[2751:2736];
    adder_tree_tier_1_p0_in[1391:1376] = adder_tree_tier_0_p0_in[2767:2752] + adder_tree_tier_0_p0_in[2783:2768];
    adder_tree_tier_1_p0_in[1407:1392] = adder_tree_tier_0_p0_in[2799:2784] + adder_tree_tier_0_p0_in[2815:2800];
    adder_tree_tier_1_p0_in[1423:1408] = adder_tree_tier_0_p0_in[2831:2816] + adder_tree_tier_0_p0_in[2847:2832];
    adder_tree_tier_1_p0_in[1439:1424] = adder_tree_tier_0_p0_in[2863:2848] + adder_tree_tier_0_p0_in[2879:2864];
    adder_tree_tier_1_p0_in[1455:1440] = adder_tree_tier_0_p0_in[2895:2880] + adder_tree_tier_0_p0_in[2911:2896];
    adder_tree_tier_1_p0_in[1471:1456] = adder_tree_tier_0_p0_in[2927:2912] + adder_tree_tier_0_p0_in[2943:2928];
    adder_tree_tier_1_p0_in[1487:1472] = adder_tree_tier_0_p0_in[2959:2944] + adder_tree_tier_0_p0_in[2975:2960];
    adder_tree_tier_1_p0_in[1503:1488] = adder_tree_tier_0_p0_in[2991:2976] + adder_tree_tier_0_p0_in[3007:2992];
    adder_tree_tier_1_p0_in[1519:1504] = adder_tree_tier_0_p0_in[3023:3008] + adder_tree_tier_0_p0_in[3039:3024];
    adder_tree_tier_1_p0_in[1535:1520] = adder_tree_tier_0_p0_in[3055:3040] + adder_tree_tier_0_p0_in[3071:3056];
    adder_tree_tier_1_p0_in[1551:1536] = adder_tree_tier_0_p0_in[3087:3072] + adder_tree_tier_0_p0_in[3103:3088];
    adder_tree_tier_1_p0_in[1567:1552] = adder_tree_tier_0_p0_in[3119:3104] + adder_tree_tier_0_p0_in[3135:3120];
    adder_tree_tier_1_p0_in[1583:1568] = adder_tree_tier_0_p0_in[3151:3136] + adder_tree_tier_0_p0_in[3167:3152];
    adder_tree_tier_1_p0_in[1599:1584] = adder_tree_tier_0_p0_in[3183:3168] + adder_tree_tier_0_p0_in[3199:3184];
    adder_tree_tier_1_p0_in[1615:1600] = adder_tree_tier_0_p0_in[3215:3200] + adder_tree_tier_0_p0_in[3231:3216];
    adder_tree_tier_1_p0_in[1631:1616] = adder_tree_tier_0_p0_in[3247:3232] + adder_tree_tier_0_p0_in[3263:3248];
    adder_tree_tier_1_p0_in[1647:1632] = adder_tree_tier_0_p0_in[3279:3264] + adder_tree_tier_0_p0_in[3295:3280];
    adder_tree_tier_1_p0_in[1663:1648] = adder_tree_tier_0_p0_in[3311:3296] + adder_tree_tier_0_p0_in[3327:3312];
    adder_tree_tier_1_p0_in[1679:1664] = adder_tree_tier_0_p0_in[3343:3328] + adder_tree_tier_0_p0_in[3359:3344];
    adder_tree_tier_1_p0_in[1695:1680] = adder_tree_tier_0_p0_in[3375:3360] + adder_tree_tier_0_p0_in[3391:3376];
    adder_tree_tier_1_p0_in[1711:1696] = adder_tree_tier_0_p0_in[3407:3392] + adder_tree_tier_0_p0_in[3423:3408];
    adder_tree_tier_1_p0_in[1727:1712] = adder_tree_tier_0_p0_in[3439:3424] + adder_tree_tier_0_p0_in[3455:3440];
    adder_tree_tier_1_p0_in[1743:1728] = adder_tree_tier_0_p0_in[3471:3456] + adder_tree_tier_0_p0_in[3487:3472];
    adder_tree_tier_1_p0_in[1759:1744] = adder_tree_tier_0_p0_in[3503:3488] + adder_tree_tier_0_p0_in[3519:3504];
    adder_tree_tier_1_p0_in[1775:1760] = adder_tree_tier_0_p0_in[3535:3520] + adder_tree_tier_0_p0_in[3551:3536];
    adder_tree_tier_1_p0_in[1791:1776] = adder_tree_tier_0_p0_in[3567:3552] + adder_tree_tier_0_p0_in[3583:3568];
    adder_tree_tier_1_p0_in[1807:1792] = adder_tree_tier_0_p0_in[3599:3584] + adder_tree_tier_0_p0_in[3615:3600];
    adder_tree_tier_1_p0_in[1823:1808] = adder_tree_tier_0_p0_in[3631:3616] + adder_tree_tier_0_p0_in[3647:3632];
    adder_tree_tier_1_p0_in[1839:1824] = adder_tree_tier_0_p0_in[3663:3648] + adder_tree_tier_0_p0_in[3679:3664];
    adder_tree_tier_1_p0_in[1855:1840] = adder_tree_tier_0_p0_in[3695:3680] + adder_tree_tier_0_p0_in[3711:3696];
    adder_tree_tier_1_p0_in[1871:1856] = adder_tree_tier_0_p0_in[3727:3712] + adder_tree_tier_0_p0_in[3743:3728];
    adder_tree_tier_1_p0_in[1887:1872] = adder_tree_tier_0_p0_in[3759:3744] + adder_tree_tier_0_p0_in[3775:3760];
    adder_tree_tier_1_p0_in[1903:1888] = adder_tree_tier_0_p0_in[3791:3776] + adder_tree_tier_0_p0_in[3807:3792];
    adder_tree_tier_1_p0_in[1919:1904] = adder_tree_tier_0_p0_in[3823:3808] + adder_tree_tier_0_p0_in[3839:3824];
    adder_tree_tier_1_p0_in[1935:1920] = adder_tree_tier_0_p0_in[3855:3840] + adder_tree_tier_0_p0_in[3871:3856];
    adder_tree_tier_1_p0_in[1951:1936] = adder_tree_tier_0_p0_in[3887:3872] + adder_tree_tier_0_p0_in[3903:3888];
    adder_tree_tier_1_p0_in[1967:1952] = adder_tree_tier_0_p0_in[3919:3904] + adder_tree_tier_0_p0_in[3935:3920];
    adder_tree_tier_1_p0_in[1983:1968] = adder_tree_tier_0_p0_in[3951:3936] + adder_tree_tier_0_p0_in[3967:3952];
    adder_tree_tier_1_p0_in[1999:1984] = adder_tree_tier_0_p0_in[3983:3968] + adder_tree_tier_0_p0_in[3999:3984];
    adder_tree_tier_1_p0_in[2015:2000] = adder_tree_tier_0_p0_in[4015:4000] + adder_tree_tier_0_p0_in[4031:4016];
    adder_tree_tier_1_p0_in[2031:2016] = adder_tree_tier_0_p0_in[4047:4032] + adder_tree_tier_0_p0_in[4063:4048];
    adder_tree_tier_1_p0_in[2047:2032] = adder_tree_tier_0_p0_in[4079:4064] + adder_tree_tier_0_p0_in[4095:4080];
    adder_tree_tier_1_p0_in[2063:2048] = adder_tree_tier_0_p0_in[4111:4096] + adder_tree_tier_0_p0_in[4127:4112];
    adder_tree_tier_1_p0_in[2079:2064] = adder_tree_tier_0_p0_in[4143:4128] + adder_tree_tier_0_p0_in[4159:4144];
    adder_tree_tier_1_p0_in[2095:2080] = adder_tree_tier_0_p0_in[4175:4160] + adder_tree_tier_0_p0_in[4191:4176];
    adder_tree_tier_1_p0_in[2111:2096] = adder_tree_tier_0_p0_in[4207:4192] + adder_tree_tier_0_p0_in[4223:4208];
    adder_tree_tier_1_p0_in[2127:2112] = adder_tree_tier_0_p0_in[4239:4224] + adder_tree_tier_0_p0_in[4255:4240];
    adder_tree_tier_1_p0_in[2143:2128] = adder_tree_tier_0_p0_in[4271:4256] + adder_tree_tier_0_p0_in[4287:4272];
    adder_tree_tier_1_p0_in[2159:2144] = adder_tree_tier_0_p0_in[4303:4288] + adder_tree_tier_0_p0_in[4319:4304];
    adder_tree_tier_1_p0_in[2175:2160] = adder_tree_tier_0_p0_in[4335:4320] + adder_tree_tier_0_p0_in[4351:4336];
    adder_tree_tier_1_p0_in[2191:2176] = adder_tree_tier_0_p0_in[4367:4352] + adder_tree_tier_0_p0_in[4383:4368];
    adder_tree_tier_1_p0_in[2207:2192] = adder_tree_tier_0_p0_in[4399:4384] + adder_tree_tier_0_p0_in[4415:4400];
    adder_tree_tier_1_p0_in[2223:2208] = adder_tree_tier_0_p0_in[4431:4416] + adder_tree_tier_0_p0_in[4447:4432];
    adder_tree_tier_1_p0_in[2239:2224] = adder_tree_tier_0_p0_in[4463:4448] + adder_tree_tier_0_p0_in[4479:4464];
    adder_tree_tier_1_p0_in[2255:2240] = adder_tree_tier_0_p0_in[4495:4480] + adder_tree_tier_0_p0_in[4511:4496];
    adder_tree_tier_1_p0_in[2271:2256] = adder_tree_tier_0_p0_in[4527:4512] + adder_tree_tier_0_p0_in[4543:4528];
    adder_tree_tier_1_p0_in[2287:2272] = adder_tree_tier_0_p0_in[4559:4544] + adder_tree_tier_0_p0_in[4575:4560];
    adder_tree_tier_1_p0_in[2303:2288] = adder_tree_tier_0_p0_in[4591:4576] + adder_tree_tier_0_p0_in[4607:4592];
    adder_tree_tier_1_p0_in[2319:2304] = adder_tree_tier_0_p0_in[4623:4608] + adder_tree_tier_0_p0_in[4639:4624];
    adder_tree_tier_1_p0_in[2335:2320] = adder_tree_tier_0_p0_in[4655:4640] + adder_tree_tier_0_p0_in[4671:4656];
    adder_tree_tier_1_p0_in[2351:2336] = adder_tree_tier_0_p0_in[4687:4672] + adder_tree_tier_0_p0_in[4703:4688];
    adder_tree_tier_1_p0_in[2367:2352] = adder_tree_tier_0_p0_in[4719:4704] + adder_tree_tier_0_p0_in[4735:4720];
    adder_tree_tier_1_p0_in[2383:2368] = adder_tree_tier_0_p0_in[4751:4736] + adder_tree_tier_0_p0_in[4767:4752];
    adder_tree_tier_1_p0_in[2399:2384] = adder_tree_tier_0_p0_in[4783:4768] + adder_tree_tier_0_p0_in[4799:4784];
    adder_tree_tier_1_p0_in[2415:2400] = adder_tree_tier_0_p0_in[4815:4800] + adder_tree_tier_0_p0_in[4831:4816];
    adder_tree_tier_1_p0_in[2431:2416] = adder_tree_tier_0_p0_in[4847:4832] + adder_tree_tier_0_p0_in[4863:4848];
    adder_tree_tier_1_p0_in[2447:2432] = adder_tree_tier_0_p0_in[4879:4864] + adder_tree_tier_0_p0_in[4895:4880];
    adder_tree_tier_1_p0_in[2463:2448] = adder_tree_tier_0_p0_in[4911:4896] + adder_tree_tier_0_p0_in[4927:4912];
    adder_tree_tier_1_p0_in[2479:2464] = adder_tree_tier_0_p0_in[4943:4928] + adder_tree_tier_0_p0_in[4959:4944];
    adder_tree_tier_1_p0_in[2495:2480] = adder_tree_tier_0_p0_in[4975:4960] + adder_tree_tier_0_p0_in[4991:4976];
    adder_tree_tier_1_p0_in[2511:2496] = adder_tree_tier_0_p0_in[5007:4992] + adder_tree_tier_0_p0_in[5023:5008];
    adder_tree_tier_1_p0_in[2527:2512] = adder_tree_tier_0_p0_in[5039:5024] + adder_tree_tier_0_p0_in[5055:5040];
    adder_tree_tier_1_p0_in[2543:2528] = adder_tree_tier_0_p0_in[5071:5056] + adder_tree_tier_0_p0_in[5087:5072];
    adder_tree_tier_1_p0_in[2559:2544] = adder_tree_tier_0_p0_in[5103:5088] + adder_tree_tier_0_p0_in[5119:5104];
    adder_tree_tier_1_p0_in[2575:2560] = adder_tree_tier_0_p0_in[5135:5120] + adder_tree_tier_0_p0_in[5151:5136];
    adder_tree_tier_1_p0_in[2591:2576] = adder_tree_tier_0_p0_in[5167:5152] + adder_tree_tier_0_p0_in[5183:5168];
    adder_tree_tier_1_p0_in[2607:2592] = adder_tree_tier_0_p0_in[5199:5184] + adder_tree_tier_0_p0_in[5215:5200];
    adder_tree_tier_1_p0_in[2623:2608] = adder_tree_tier_0_p0_in[5231:5216] + adder_tree_tier_0_p0_in[5247:5232];
    adder_tree_tier_1_p0_in[2639:2624] = adder_tree_tier_0_p0_in[5263:5248] + adder_tree_tier_0_p0_in[5279:5264];
    adder_tree_tier_1_p0_in[2655:2640] = adder_tree_tier_0_p0_in[5295:5280] + adder_tree_tier_0_p0_in[5311:5296];
    adder_tree_tier_1_p0_in[2671:2656] = adder_tree_tier_0_p0_in[5327:5312] + adder_tree_tier_0_p0_in[5343:5328];
    adder_tree_tier_1_p0_in[2687:2672] = adder_tree_tier_0_p0_in[5359:5344] + adder_tree_tier_0_p0_in[5375:5360];
    adder_tree_tier_1_p0_in[2703:2688] = adder_tree_tier_0_p0_in[5391:5376] + adder_tree_tier_0_p0_in[5407:5392];
    adder_tree_tier_1_p0_in[2719:2704] = adder_tree_tier_0_p0_in[5423:5408] + adder_tree_tier_0_p0_in[5439:5424];
    adder_tree_tier_1_p0_in[2735:2720] = adder_tree_tier_0_p0_in[5455:5440] + adder_tree_tier_0_p0_in[5471:5456];
    adder_tree_tier_1_p0_in[2751:2736] = adder_tree_tier_0_p0_in[5487:5472] + adder_tree_tier_0_p0_in[5503:5488];
    adder_tree_tier_1_p0_in[2767:2752] = adder_tree_tier_0_p0_in[5519:5504] + adder_tree_tier_0_p0_in[5535:5520];
    adder_tree_tier_1_p0_in[2783:2768] = adder_tree_tier_0_p0_in[5551:5536] + adder_tree_tier_0_p0_in[5567:5552];
    adder_tree_tier_1_p0_in[2799:2784] = adder_tree_tier_0_p0_in[5583:5568] + adder_tree_tier_0_p0_in[5599:5584];
    adder_tree_tier_1_p0_in[2815:2800] = adder_tree_tier_0_p0_in[5615:5600] + adder_tree_tier_0_p0_in[5631:5616];
    adder_tree_tier_1_p0_in[2831:2816] = adder_tree_tier_0_p0_in[5647:5632] + adder_tree_tier_0_p0_in[5663:5648];
    adder_tree_tier_1_p0_in[2847:2832] = adder_tree_tier_0_p0_in[5679:5664] + adder_tree_tier_0_p0_in[5695:5680];
    adder_tree_tier_1_p0_in[2863:2848] = adder_tree_tier_0_p0_in[5711:5696] + adder_tree_tier_0_p0_in[5727:5712];
    adder_tree_tier_1_p0_in[2879:2864] = adder_tree_tier_0_p0_in[5743:5728] + adder_tree_tier_0_p0_in[5759:5744];
    adder_tree_tier_1_p0_in[2895:2880] = adder_tree_tier_0_p0_in[5775:5760] + adder_tree_tier_0_p0_in[5791:5776];
    adder_tree_tier_1_p0_in[2911:2896] = adder_tree_tier_0_p0_in[5807:5792] + adder_tree_tier_0_p0_in[5823:5808];
    adder_tree_tier_1_p0_in[2927:2912] = adder_tree_tier_0_p0_in[5839:5824] + adder_tree_tier_0_p0_in[5855:5840];
    adder_tree_tier_1_p0_in[2943:2928] = adder_tree_tier_0_p0_in[5871:5856] + adder_tree_tier_0_p0_in[5887:5872];
    adder_tree_tier_1_p0_in[2959:2944] = adder_tree_tier_0_p0_in[5903:5888] + adder_tree_tier_0_p0_in[5919:5904];
    adder_tree_tier_1_p0_in[2975:2960] = adder_tree_tier_0_p0_in[5935:5920] + adder_tree_tier_0_p0_in[5951:5936];
    adder_tree_tier_1_p0_in[2991:2976] = adder_tree_tier_0_p0_in[5967:5952] + adder_tree_tier_0_p0_in[5983:5968];
    adder_tree_tier_1_p0_in[3007:2992] = adder_tree_tier_0_p0_in[5999:5984] + adder_tree_tier_0_p0_in[6015:6000];
    adder_tree_tier_1_p0_in[3023:3008] = adder_tree_tier_0_p0_in[6031:6016] + adder_tree_tier_0_p0_in[6047:6032];
    adder_tree_tier_1_p0_in[3039:3024] = adder_tree_tier_0_p0_in[6063:6048] + adder_tree_tier_0_p0_in[6079:6064];
    adder_tree_tier_1_p0_in[3055:3040] = adder_tree_tier_0_p0_in[6095:6080] + adder_tree_tier_0_p0_in[6111:6096];
    adder_tree_tier_1_p0_in[3071:3056] = adder_tree_tier_0_p0_in[6127:6112] + adder_tree_tier_0_p0_in[6143:6128];
    adder_tree_tier_1_p0_in[3087:3072] = adder_tree_tier_0_p0_in[6159:6144] + adder_tree_tier_0_p0_in[6175:6160];
    adder_tree_tier_1_p0_in[3103:3088] = adder_tree_tier_0_p0_in[6191:6176] + adder_tree_tier_0_p0_in[6207:6192];
    adder_tree_tier_1_p0_in[3119:3104] = adder_tree_tier_0_p0_in[6223:6208] + adder_tree_tier_0_p0_in[6239:6224];
    adder_tree_tier_1_p0_in[3135:3120] = adder_tree_tier_0_p0_in[6255:6240] + adder_tree_tier_0_p0_in[6271:6256];
    adder_tree_tier_1_p0_in[3151:3136] = adder_tree_tier_0_p0_in[6287:6272] + adder_tree_tier_0_p0_in[6303:6288];
    adder_tree_tier_1_p0_in[3167:3152] = adder_tree_tier_0_p0_in[6319:6304] + adder_tree_tier_0_p0_in[6335:6320];
    adder_tree_tier_1_p0_in[3183:3168] = adder_tree_tier_0_p0_in[6351:6336] + adder_tree_tier_0_p0_in[6367:6352];
    adder_tree_tier_1_p0_in[3199:3184] = adder_tree_tier_0_p0_in[6383:6368] + adder_tree_tier_0_p0_in[6399:6384];
    adder_tree_tier_1_p0_in[3215:3200] = adder_tree_tier_0_p0_in[6415:6400];
    adder_tree_tier_2_p0_in[15:0] = adder_tree_tier_1_p0_in[15:0] + adder_tree_tier_1_p0_in[31:16];
    adder_tree_tier_2_p0_in[31:16] = adder_tree_tier_1_p0_in[47:32] + adder_tree_tier_1_p0_in[63:48];
    adder_tree_tier_2_p0_in[47:32] = adder_tree_tier_1_p0_in[79:64] + adder_tree_tier_1_p0_in[95:80];
    adder_tree_tier_2_p0_in[63:48] = adder_tree_tier_1_p0_in[111:96] + adder_tree_tier_1_p0_in[127:112];
    adder_tree_tier_2_p0_in[79:64] = adder_tree_tier_1_p0_in[143:128] + adder_tree_tier_1_p0_in[159:144];
    adder_tree_tier_2_p0_in[95:80] = adder_tree_tier_1_p0_in[175:160] + adder_tree_tier_1_p0_in[191:176];
    adder_tree_tier_2_p0_in[111:96] = adder_tree_tier_1_p0_in[207:192] + adder_tree_tier_1_p0_in[223:208];
    adder_tree_tier_2_p0_in[127:112] = adder_tree_tier_1_p0_in[239:224] + adder_tree_tier_1_p0_in[255:240];
    adder_tree_tier_2_p0_in[143:128] = adder_tree_tier_1_p0_in[271:256] + adder_tree_tier_1_p0_in[287:272];
    adder_tree_tier_2_p0_in[159:144] = adder_tree_tier_1_p0_in[303:288] + adder_tree_tier_1_p0_in[319:304];
    adder_tree_tier_2_p0_in[175:160] = adder_tree_tier_1_p0_in[335:320] + adder_tree_tier_1_p0_in[351:336];
    adder_tree_tier_2_p0_in[191:176] = adder_tree_tier_1_p0_in[367:352] + adder_tree_tier_1_p0_in[383:368];
    adder_tree_tier_2_p0_in[207:192] = adder_tree_tier_1_p0_in[399:384] + adder_tree_tier_1_p0_in[415:400];
    adder_tree_tier_2_p0_in[223:208] = adder_tree_tier_1_p0_in[431:416] + adder_tree_tier_1_p0_in[447:432];
    adder_tree_tier_2_p0_in[239:224] = adder_tree_tier_1_p0_in[463:448] + adder_tree_tier_1_p0_in[479:464];
    adder_tree_tier_2_p0_in[255:240] = adder_tree_tier_1_p0_in[495:480] + adder_tree_tier_1_p0_in[511:496];
    adder_tree_tier_2_p0_in[271:256] = adder_tree_tier_1_p0_in[527:512] + adder_tree_tier_1_p0_in[543:528];
    adder_tree_tier_2_p0_in[287:272] = adder_tree_tier_1_p0_in[559:544] + adder_tree_tier_1_p0_in[575:560];
    adder_tree_tier_2_p0_in[303:288] = adder_tree_tier_1_p0_in[591:576] + adder_tree_tier_1_p0_in[607:592];
    adder_tree_tier_2_p0_in[319:304] = adder_tree_tier_1_p0_in[623:608] + adder_tree_tier_1_p0_in[639:624];
    adder_tree_tier_2_p0_in[335:320] = adder_tree_tier_1_p0_in[655:640] + adder_tree_tier_1_p0_in[671:656];
    adder_tree_tier_2_p0_in[351:336] = adder_tree_tier_1_p0_in[687:672] + adder_tree_tier_1_p0_in[703:688];
    adder_tree_tier_2_p0_in[367:352] = adder_tree_tier_1_p0_in[719:704] + adder_tree_tier_1_p0_in[735:720];
    adder_tree_tier_2_p0_in[383:368] = adder_tree_tier_1_p0_in[751:736] + adder_tree_tier_1_p0_in[767:752];
    adder_tree_tier_2_p0_in[399:384] = adder_tree_tier_1_p0_in[783:768] + adder_tree_tier_1_p0_in[799:784];
    adder_tree_tier_2_p0_in[415:400] = adder_tree_tier_1_p0_in[815:800] + adder_tree_tier_1_p0_in[831:816];
    adder_tree_tier_2_p0_in[431:416] = adder_tree_tier_1_p0_in[847:832] + adder_tree_tier_1_p0_in[863:848];
    adder_tree_tier_2_p0_in[447:432] = adder_tree_tier_1_p0_in[879:864] + adder_tree_tier_1_p0_in[895:880];
    adder_tree_tier_2_p0_in[463:448] = adder_tree_tier_1_p0_in[911:896] + adder_tree_tier_1_p0_in[927:912];
    adder_tree_tier_2_p0_in[479:464] = adder_tree_tier_1_p0_in[943:928] + adder_tree_tier_1_p0_in[959:944];
    adder_tree_tier_2_p0_in[495:480] = adder_tree_tier_1_p0_in[975:960] + adder_tree_tier_1_p0_in[991:976];
    adder_tree_tier_2_p0_in[511:496] = adder_tree_tier_1_p0_in[1007:992] + adder_tree_tier_1_p0_in[1023:1008];
    adder_tree_tier_2_p0_in[527:512] = adder_tree_tier_1_p0_in[1039:1024] + adder_tree_tier_1_p0_in[1055:1040];
    adder_tree_tier_2_p0_in[543:528] = adder_tree_tier_1_p0_in[1071:1056] + adder_tree_tier_1_p0_in[1087:1072];
    adder_tree_tier_2_p0_in[559:544] = adder_tree_tier_1_p0_in[1103:1088] + adder_tree_tier_1_p0_in[1119:1104];
    adder_tree_tier_2_p0_in[575:560] = adder_tree_tier_1_p0_in[1135:1120] + adder_tree_tier_1_p0_in[1151:1136];
    adder_tree_tier_2_p0_in[591:576] = adder_tree_tier_1_p0_in[1167:1152] + adder_tree_tier_1_p0_in[1183:1168];
    adder_tree_tier_2_p0_in[607:592] = adder_tree_tier_1_p0_in[1199:1184] + adder_tree_tier_1_p0_in[1215:1200];
    adder_tree_tier_2_p0_in[623:608] = adder_tree_tier_1_p0_in[1231:1216] + adder_tree_tier_1_p0_in[1247:1232];
    adder_tree_tier_2_p0_in[639:624] = adder_tree_tier_1_p0_in[1263:1248] + adder_tree_tier_1_p0_in[1279:1264];
    adder_tree_tier_2_p0_in[655:640] = adder_tree_tier_1_p0_in[1295:1280] + adder_tree_tier_1_p0_in[1311:1296];
    adder_tree_tier_2_p0_in[671:656] = adder_tree_tier_1_p0_in[1327:1312] + adder_tree_tier_1_p0_in[1343:1328];
    adder_tree_tier_2_p0_in[687:672] = adder_tree_tier_1_p0_in[1359:1344] + adder_tree_tier_1_p0_in[1375:1360];
    adder_tree_tier_2_p0_in[703:688] = adder_tree_tier_1_p0_in[1391:1376] + adder_tree_tier_1_p0_in[1407:1392];
    adder_tree_tier_2_p0_in[719:704] = adder_tree_tier_1_p0_in[1423:1408] + adder_tree_tier_1_p0_in[1439:1424];
    adder_tree_tier_2_p0_in[735:720] = adder_tree_tier_1_p0_in[1455:1440] + adder_tree_tier_1_p0_in[1471:1456];
    adder_tree_tier_2_p0_in[751:736] = adder_tree_tier_1_p0_in[1487:1472] + adder_tree_tier_1_p0_in[1503:1488];
    adder_tree_tier_2_p0_in[767:752] = adder_tree_tier_1_p0_in[1519:1504] + adder_tree_tier_1_p0_in[1535:1520];
    adder_tree_tier_2_p0_in[783:768] = adder_tree_tier_1_p0_in[1551:1536] + adder_tree_tier_1_p0_in[1567:1552];
    adder_tree_tier_2_p0_in[799:784] = adder_tree_tier_1_p0_in[1583:1568] + adder_tree_tier_1_p0_in[1599:1584];
    adder_tree_tier_2_p0_in[815:800] = adder_tree_tier_1_p0_in[1615:1600] + adder_tree_tier_1_p0_in[1631:1616];
    adder_tree_tier_2_p0_in[831:816] = adder_tree_tier_1_p0_in[1647:1632] + adder_tree_tier_1_p0_in[1663:1648];
    adder_tree_tier_2_p0_in[847:832] = adder_tree_tier_1_p0_in[1679:1664] + adder_tree_tier_1_p0_in[1695:1680];
    adder_tree_tier_2_p0_in[863:848] = adder_tree_tier_1_p0_in[1711:1696] + adder_tree_tier_1_p0_in[1727:1712];
    adder_tree_tier_2_p0_in[879:864] = adder_tree_tier_1_p0_in[1743:1728] + adder_tree_tier_1_p0_in[1759:1744];
    adder_tree_tier_2_p0_in[895:880] = adder_tree_tier_1_p0_in[1775:1760] + adder_tree_tier_1_p0_in[1791:1776];
    adder_tree_tier_2_p0_in[911:896] = adder_tree_tier_1_p0_in[1807:1792] + adder_tree_tier_1_p0_in[1823:1808];
    adder_tree_tier_2_p0_in[927:912] = adder_tree_tier_1_p0_in[1839:1824] + adder_tree_tier_1_p0_in[1855:1840];
    adder_tree_tier_2_p0_in[943:928] = adder_tree_tier_1_p0_in[1871:1856] + adder_tree_tier_1_p0_in[1887:1872];
    adder_tree_tier_2_p0_in[959:944] = adder_tree_tier_1_p0_in[1903:1888] + adder_tree_tier_1_p0_in[1919:1904];
    adder_tree_tier_2_p0_in[975:960] = adder_tree_tier_1_p0_in[1935:1920] + adder_tree_tier_1_p0_in[1951:1936];
    adder_tree_tier_2_p0_in[991:976] = adder_tree_tier_1_p0_in[1967:1952] + adder_tree_tier_1_p0_in[1983:1968];
    adder_tree_tier_2_p0_in[1007:992] = adder_tree_tier_1_p0_in[1999:1984] + adder_tree_tier_1_p0_in[2015:2000];
    adder_tree_tier_2_p0_in[1023:1008] = adder_tree_tier_1_p0_in[2031:2016] + adder_tree_tier_1_p0_in[2047:2032];
    adder_tree_tier_2_p0_in[1039:1024] = adder_tree_tier_1_p0_in[2063:2048] + adder_tree_tier_1_p0_in[2079:2064];
    adder_tree_tier_2_p0_in[1055:1040] = adder_tree_tier_1_p0_in[2095:2080] + adder_tree_tier_1_p0_in[2111:2096];
    adder_tree_tier_2_p0_in[1071:1056] = adder_tree_tier_1_p0_in[2127:2112] + adder_tree_tier_1_p0_in[2143:2128];
    adder_tree_tier_2_p0_in[1087:1072] = adder_tree_tier_1_p0_in[2159:2144] + adder_tree_tier_1_p0_in[2175:2160];
    adder_tree_tier_2_p0_in[1103:1088] = adder_tree_tier_1_p0_in[2191:2176] + adder_tree_tier_1_p0_in[2207:2192];
    adder_tree_tier_2_p0_in[1119:1104] = adder_tree_tier_1_p0_in[2223:2208] + adder_tree_tier_1_p0_in[2239:2224];
    adder_tree_tier_2_p0_in[1135:1120] = adder_tree_tier_1_p0_in[2255:2240] + adder_tree_tier_1_p0_in[2271:2256];
    adder_tree_tier_2_p0_in[1151:1136] = adder_tree_tier_1_p0_in[2287:2272] + adder_tree_tier_1_p0_in[2303:2288];
    adder_tree_tier_2_p0_in[1167:1152] = adder_tree_tier_1_p0_in[2319:2304] + adder_tree_tier_1_p0_in[2335:2320];
    adder_tree_tier_2_p0_in[1183:1168] = adder_tree_tier_1_p0_in[2351:2336] + adder_tree_tier_1_p0_in[2367:2352];
    adder_tree_tier_2_p0_in[1199:1184] = adder_tree_tier_1_p0_in[2383:2368] + adder_tree_tier_1_p0_in[2399:2384];
    adder_tree_tier_2_p0_in[1215:1200] = adder_tree_tier_1_p0_in[2415:2400] + adder_tree_tier_1_p0_in[2431:2416];
    adder_tree_tier_2_p0_in[1231:1216] = adder_tree_tier_1_p0_in[2447:2432] + adder_tree_tier_1_p0_in[2463:2448];
    adder_tree_tier_2_p0_in[1247:1232] = adder_tree_tier_1_p0_in[2479:2464] + adder_tree_tier_1_p0_in[2495:2480];
    adder_tree_tier_2_p0_in[1263:1248] = adder_tree_tier_1_p0_in[2511:2496] + adder_tree_tier_1_p0_in[2527:2512];
    adder_tree_tier_2_p0_in[1279:1264] = adder_tree_tier_1_p0_in[2543:2528] + adder_tree_tier_1_p0_in[2559:2544];
    adder_tree_tier_2_p0_in[1295:1280] = adder_tree_tier_1_p0_in[2575:2560] + adder_tree_tier_1_p0_in[2591:2576];
    adder_tree_tier_2_p0_in[1311:1296] = adder_tree_tier_1_p0_in[2607:2592] + adder_tree_tier_1_p0_in[2623:2608];
    adder_tree_tier_2_p0_in[1327:1312] = adder_tree_tier_1_p0_in[2639:2624] + adder_tree_tier_1_p0_in[2655:2640];
    adder_tree_tier_2_p0_in[1343:1328] = adder_tree_tier_1_p0_in[2671:2656] + adder_tree_tier_1_p0_in[2687:2672];
    adder_tree_tier_2_p0_in[1359:1344] = adder_tree_tier_1_p0_in[2703:2688] + adder_tree_tier_1_p0_in[2719:2704];
    adder_tree_tier_2_p0_in[1375:1360] = adder_tree_tier_1_p0_in[2735:2720] + adder_tree_tier_1_p0_in[2751:2736];
    adder_tree_tier_2_p0_in[1391:1376] = adder_tree_tier_1_p0_in[2767:2752] + adder_tree_tier_1_p0_in[2783:2768];
    adder_tree_tier_2_p0_in[1407:1392] = adder_tree_tier_1_p0_in[2799:2784] + adder_tree_tier_1_p0_in[2815:2800];
    adder_tree_tier_2_p0_in[1423:1408] = adder_tree_tier_1_p0_in[2831:2816] + adder_tree_tier_1_p0_in[2847:2832];
    adder_tree_tier_2_p0_in[1439:1424] = adder_tree_tier_1_p0_in[2863:2848] + adder_tree_tier_1_p0_in[2879:2864];
    adder_tree_tier_2_p0_in[1455:1440] = adder_tree_tier_1_p0_in[2895:2880] + adder_tree_tier_1_p0_in[2911:2896];
    adder_tree_tier_2_p0_in[1471:1456] = adder_tree_tier_1_p0_in[2927:2912] + adder_tree_tier_1_p0_in[2943:2928];
    adder_tree_tier_2_p0_in[1487:1472] = adder_tree_tier_1_p0_in[2959:2944] + adder_tree_tier_1_p0_in[2975:2960];
    adder_tree_tier_2_p0_in[1503:1488] = adder_tree_tier_1_p0_in[2991:2976] + adder_tree_tier_1_p0_in[3007:2992];
    adder_tree_tier_2_p0_in[1519:1504] = adder_tree_tier_1_p0_in[3023:3008] + adder_tree_tier_1_p0_in[3039:3024];
    adder_tree_tier_2_p0_in[1535:1520] = adder_tree_tier_1_p0_in[3055:3040] + adder_tree_tier_1_p0_in[3071:3056];
    adder_tree_tier_2_p0_in[1551:1536] = adder_tree_tier_1_p0_in[3087:3072] + adder_tree_tier_1_p0_in[3103:3088];
    adder_tree_tier_2_p0_in[1567:1552] = adder_tree_tier_1_p0_in[3119:3104] + adder_tree_tier_1_p0_in[3135:3120];
    adder_tree_tier_2_p0_in[1583:1568] = adder_tree_tier_1_p0_in[3151:3136] + adder_tree_tier_1_p0_in[3167:3152];
    adder_tree_tier_2_p0_in[1599:1584] = adder_tree_tier_1_p0_in[3183:3168] + adder_tree_tier_1_p0_in[3199:3184];
    adder_tree_tier_2_p0_in[1615:1600] = adder_tree_tier_1_p0_in[3215:3200];
    adder_tree_tier_3_p0_in[15:0] = adder_tree_tier_2_p0_in[15:0] + adder_tree_tier_2_p0_in[31:16];
    adder_tree_tier_3_p0_in[31:16] = adder_tree_tier_2_p0_in[47:32] + adder_tree_tier_2_p0_in[63:48];
    adder_tree_tier_3_p0_in[47:32] = adder_tree_tier_2_p0_in[79:64] + adder_tree_tier_2_p0_in[95:80];
    adder_tree_tier_3_p0_in[63:48] = adder_tree_tier_2_p0_in[111:96] + adder_tree_tier_2_p0_in[127:112];
    adder_tree_tier_3_p0_in[79:64] = adder_tree_tier_2_p0_in[143:128] + adder_tree_tier_2_p0_in[159:144];
    adder_tree_tier_3_p0_in[95:80] = adder_tree_tier_2_p0_in[175:160] + adder_tree_tier_2_p0_in[191:176];
    adder_tree_tier_3_p0_in[111:96] = adder_tree_tier_2_p0_in[207:192] + adder_tree_tier_2_p0_in[223:208];
    adder_tree_tier_3_p0_in[127:112] = adder_tree_tier_2_p0_in[239:224] + adder_tree_tier_2_p0_in[255:240];
    adder_tree_tier_3_p0_in[143:128] = adder_tree_tier_2_p0_in[271:256] + adder_tree_tier_2_p0_in[287:272];
    adder_tree_tier_3_p0_in[159:144] = adder_tree_tier_2_p0_in[303:288] + adder_tree_tier_2_p0_in[319:304];
    adder_tree_tier_3_p0_in[175:160] = adder_tree_tier_2_p0_in[335:320] + adder_tree_tier_2_p0_in[351:336];
    adder_tree_tier_3_p0_in[191:176] = adder_tree_tier_2_p0_in[367:352] + adder_tree_tier_2_p0_in[383:368];
    adder_tree_tier_3_p0_in[207:192] = adder_tree_tier_2_p0_in[399:384] + adder_tree_tier_2_p0_in[415:400];
    adder_tree_tier_3_p0_in[223:208] = adder_tree_tier_2_p0_in[431:416] + adder_tree_tier_2_p0_in[447:432];
    adder_tree_tier_3_p0_in[239:224] = adder_tree_tier_2_p0_in[463:448] + adder_tree_tier_2_p0_in[479:464];
    adder_tree_tier_3_p0_in[255:240] = adder_tree_tier_2_p0_in[495:480] + adder_tree_tier_2_p0_in[511:496];
    adder_tree_tier_3_p0_in[271:256] = adder_tree_tier_2_p0_in[527:512] + adder_tree_tier_2_p0_in[543:528];
    adder_tree_tier_3_p0_in[287:272] = adder_tree_tier_2_p0_in[559:544] + adder_tree_tier_2_p0_in[575:560];
    adder_tree_tier_3_p0_in[303:288] = adder_tree_tier_2_p0_in[591:576] + adder_tree_tier_2_p0_in[607:592];
    adder_tree_tier_3_p0_in[319:304] = adder_tree_tier_2_p0_in[623:608] + adder_tree_tier_2_p0_in[639:624];
    adder_tree_tier_3_p0_in[335:320] = adder_tree_tier_2_p0_in[655:640] + adder_tree_tier_2_p0_in[671:656];
    adder_tree_tier_3_p0_in[351:336] = adder_tree_tier_2_p0_in[687:672] + adder_tree_tier_2_p0_in[703:688];
    adder_tree_tier_3_p0_in[367:352] = adder_tree_tier_2_p0_in[719:704] + adder_tree_tier_2_p0_in[735:720];
    adder_tree_tier_3_p0_in[383:368] = adder_tree_tier_2_p0_in[751:736] + adder_tree_tier_2_p0_in[767:752];
    adder_tree_tier_3_p0_in[399:384] = adder_tree_tier_2_p0_in[783:768] + adder_tree_tier_2_p0_in[799:784];
    adder_tree_tier_3_p0_in[415:400] = adder_tree_tier_2_p0_in[815:800] + adder_tree_tier_2_p0_in[831:816];
    adder_tree_tier_3_p0_in[431:416] = adder_tree_tier_2_p0_in[847:832] + adder_tree_tier_2_p0_in[863:848];
    adder_tree_tier_3_p0_in[447:432] = adder_tree_tier_2_p0_in[879:864] + adder_tree_tier_2_p0_in[895:880];
    adder_tree_tier_3_p0_in[463:448] = adder_tree_tier_2_p0_in[911:896] + adder_tree_tier_2_p0_in[927:912];
    adder_tree_tier_3_p0_in[479:464] = adder_tree_tier_2_p0_in[943:928] + adder_tree_tier_2_p0_in[959:944];
    adder_tree_tier_3_p0_in[495:480] = adder_tree_tier_2_p0_in[975:960] + adder_tree_tier_2_p0_in[991:976];
    adder_tree_tier_3_p0_in[511:496] = adder_tree_tier_2_p0_in[1007:992] + adder_tree_tier_2_p0_in[1023:1008];
    adder_tree_tier_3_p0_in[527:512] = adder_tree_tier_2_p0_in[1039:1024] + adder_tree_tier_2_p0_in[1055:1040];
    adder_tree_tier_3_p0_in[543:528] = adder_tree_tier_2_p0_in[1071:1056] + adder_tree_tier_2_p0_in[1087:1072];
    adder_tree_tier_3_p0_in[559:544] = adder_tree_tier_2_p0_in[1103:1088] + adder_tree_tier_2_p0_in[1119:1104];
    adder_tree_tier_3_p0_in[575:560] = adder_tree_tier_2_p0_in[1135:1120] + adder_tree_tier_2_p0_in[1151:1136];
    adder_tree_tier_3_p0_in[591:576] = adder_tree_tier_2_p0_in[1167:1152] + adder_tree_tier_2_p0_in[1183:1168];
    adder_tree_tier_3_p0_in[607:592] = adder_tree_tier_2_p0_in[1199:1184] + adder_tree_tier_2_p0_in[1215:1200];
    adder_tree_tier_3_p0_in[623:608] = adder_tree_tier_2_p0_in[1231:1216] + adder_tree_tier_2_p0_in[1247:1232];
    adder_tree_tier_3_p0_in[639:624] = adder_tree_tier_2_p0_in[1263:1248] + adder_tree_tier_2_p0_in[1279:1264];
    adder_tree_tier_3_p0_in[655:640] = adder_tree_tier_2_p0_in[1295:1280] + adder_tree_tier_2_p0_in[1311:1296];
    adder_tree_tier_3_p0_in[671:656] = adder_tree_tier_2_p0_in[1327:1312] + adder_tree_tier_2_p0_in[1343:1328];
    adder_tree_tier_3_p0_in[687:672] = adder_tree_tier_2_p0_in[1359:1344] + adder_tree_tier_2_p0_in[1375:1360];
    adder_tree_tier_3_p0_in[703:688] = adder_tree_tier_2_p0_in[1391:1376] + adder_tree_tier_2_p0_in[1407:1392];
    adder_tree_tier_3_p0_in[719:704] = adder_tree_tier_2_p0_in[1423:1408] + adder_tree_tier_2_p0_in[1439:1424];
    adder_tree_tier_3_p0_in[735:720] = adder_tree_tier_2_p0_in[1455:1440] + adder_tree_tier_2_p0_in[1471:1456];
    adder_tree_tier_3_p0_in[751:736] = adder_tree_tier_2_p0_in[1487:1472] + adder_tree_tier_2_p0_in[1503:1488];
    adder_tree_tier_3_p0_in[767:752] = adder_tree_tier_2_p0_in[1519:1504] + adder_tree_tier_2_p0_in[1535:1520];
    adder_tree_tier_3_p0_in[783:768] = adder_tree_tier_2_p0_in[1551:1536] + adder_tree_tier_2_p0_in[1567:1552];
    adder_tree_tier_3_p0_in[799:784] = adder_tree_tier_2_p0_in[1583:1568] + adder_tree_tier_2_p0_in[1599:1584];
    adder_tree_tier_3_p0_in[815:800] = adder_tree_tier_2_p0_in[1615:1600];
    adder_tree_tier_4_p0_in[15:0] = adder_tree_tier_3_p0_in[15:0] + adder_tree_tier_3_p0_in[31:16];
    adder_tree_tier_4_p0_in[31:16] = adder_tree_tier_3_p0_in[47:32] + adder_tree_tier_3_p0_in[63:48];
    adder_tree_tier_4_p0_in[47:32] = adder_tree_tier_3_p0_in[79:64] + adder_tree_tier_3_p0_in[95:80];
    adder_tree_tier_4_p0_in[63:48] = adder_tree_tier_3_p0_in[111:96] + adder_tree_tier_3_p0_in[127:112];
    adder_tree_tier_4_p0_in[79:64] = adder_tree_tier_3_p0_in[143:128] + adder_tree_tier_3_p0_in[159:144];
    adder_tree_tier_4_p0_in[95:80] = adder_tree_tier_3_p0_in[175:160] + adder_tree_tier_3_p0_in[191:176];
    adder_tree_tier_4_p0_in[111:96] = adder_tree_tier_3_p0_in[207:192] + adder_tree_tier_3_p0_in[223:208];
    adder_tree_tier_4_p0_in[127:112] = adder_tree_tier_3_p0_in[239:224] + adder_tree_tier_3_p0_in[255:240];
    adder_tree_tier_4_p0_in[143:128] = adder_tree_tier_3_p0_in[271:256] + adder_tree_tier_3_p0_in[287:272];
    adder_tree_tier_4_p0_in[159:144] = adder_tree_tier_3_p0_in[303:288] + adder_tree_tier_3_p0_in[319:304];
    adder_tree_tier_4_p0_in[175:160] = adder_tree_tier_3_p0_in[335:320] + adder_tree_tier_3_p0_in[351:336];
    adder_tree_tier_4_p0_in[191:176] = adder_tree_tier_3_p0_in[367:352] + adder_tree_tier_3_p0_in[383:368];
    adder_tree_tier_4_p0_in[207:192] = adder_tree_tier_3_p0_in[399:384] + adder_tree_tier_3_p0_in[415:400];
    adder_tree_tier_4_p0_in[223:208] = adder_tree_tier_3_p0_in[431:416] + adder_tree_tier_3_p0_in[447:432];
    adder_tree_tier_4_p0_in[239:224] = adder_tree_tier_3_p0_in[463:448] + adder_tree_tier_3_p0_in[479:464];
    adder_tree_tier_4_p0_in[255:240] = adder_tree_tier_3_p0_in[495:480] + adder_tree_tier_3_p0_in[511:496];
    adder_tree_tier_4_p0_in[271:256] = adder_tree_tier_3_p0_in[527:512] + adder_tree_tier_3_p0_in[543:528];
    adder_tree_tier_4_p0_in[287:272] = adder_tree_tier_3_p0_in[559:544] + adder_tree_tier_3_p0_in[575:560];
    adder_tree_tier_4_p0_in[303:288] = adder_tree_tier_3_p0_in[591:576] + adder_tree_tier_3_p0_in[607:592];
    adder_tree_tier_4_p0_in[319:304] = adder_tree_tier_3_p0_in[623:608] + adder_tree_tier_3_p0_in[639:624];
    adder_tree_tier_4_p0_in[335:320] = adder_tree_tier_3_p0_in[655:640] + adder_tree_tier_3_p0_in[671:656];
    adder_tree_tier_4_p0_in[351:336] = adder_tree_tier_3_p0_in[687:672] + adder_tree_tier_3_p0_in[703:688];
    adder_tree_tier_4_p0_in[367:352] = adder_tree_tier_3_p0_in[719:704] + adder_tree_tier_3_p0_in[735:720];
    adder_tree_tier_4_p0_in[383:368] = adder_tree_tier_3_p0_in[751:736] + adder_tree_tier_3_p0_in[767:752];
    adder_tree_tier_4_p0_in[399:384] = adder_tree_tier_3_p0_in[783:768] + adder_tree_tier_3_p0_in[799:784];
    adder_tree_tier_4_p0_in[415:400] = adder_tree_tier_3_p0_in[815:800];
    adder_tree_tier_5_p0_in[15:0] = adder_tree_tier_4_p0_in[15:0] + adder_tree_tier_4_p0_in[31:16];
    adder_tree_tier_5_p0_in[31:16] = adder_tree_tier_4_p0_in[47:32] + adder_tree_tier_4_p0_in[63:48];
    adder_tree_tier_5_p0_in[47:32] = adder_tree_tier_4_p0_in[79:64] + adder_tree_tier_4_p0_in[95:80];
    adder_tree_tier_5_p0_in[63:48] = adder_tree_tier_4_p0_in[111:96] + adder_tree_tier_4_p0_in[127:112];
    adder_tree_tier_5_p0_in[79:64] = adder_tree_tier_4_p0_in[143:128] + adder_tree_tier_4_p0_in[159:144];
    adder_tree_tier_5_p0_in[95:80] = adder_tree_tier_4_p0_in[175:160] + adder_tree_tier_4_p0_in[191:176];
    adder_tree_tier_5_p0_in[111:96] = adder_tree_tier_4_p0_in[207:192] + adder_tree_tier_4_p0_in[223:208];
    adder_tree_tier_5_p0_in[127:112] = adder_tree_tier_4_p0_in[239:224] + adder_tree_tier_4_p0_in[255:240];
    adder_tree_tier_5_p0_in[143:128] = adder_tree_tier_4_p0_in[271:256] + adder_tree_tier_4_p0_in[287:272];
    adder_tree_tier_5_p0_in[159:144] = adder_tree_tier_4_p0_in[303:288] + adder_tree_tier_4_p0_in[319:304];
    adder_tree_tier_5_p0_in[175:160] = adder_tree_tier_4_p0_in[335:320] + adder_tree_tier_4_p0_in[351:336];
    adder_tree_tier_5_p0_in[191:176] = adder_tree_tier_4_p0_in[367:352] + adder_tree_tier_4_p0_in[383:368];
    adder_tree_tier_5_p0_in[207:192] = adder_tree_tier_4_p0_in[399:384] + adder_tree_tier_4_p0_in[415:400];
    adder_tree_tier_6_p0_in[15:0] = adder_tree_tier_5_p0_in[15:0] + adder_tree_tier_5_p0_in[31:16];
    adder_tree_tier_6_p0_in[31:16] = adder_tree_tier_5_p0_in[47:32] + adder_tree_tier_5_p0_in[63:48];
    adder_tree_tier_6_p0_in[47:32] = adder_tree_tier_5_p0_in[79:64] + adder_tree_tier_5_p0_in[95:80];
    adder_tree_tier_6_p0_in[63:48] = adder_tree_tier_5_p0_in[111:96] + adder_tree_tier_5_p0_in[127:112];
    adder_tree_tier_6_p0_in[79:64] = adder_tree_tier_5_p0_in[143:128] + adder_tree_tier_5_p0_in[159:144];
    adder_tree_tier_6_p0_in[95:80] = adder_tree_tier_5_p0_in[175:160] + adder_tree_tier_5_p0_in[191:176];
    adder_tree_tier_6_p0_in[111:96] = adder_tree_tier_5_p0_in[207:192];
    adder_tree_tier_7_p0_in[15:0] = adder_tree_tier_6_p0_in[15:0] + adder_tree_tier_6_p0_in[31:16];
    adder_tree_tier_7_p0_in[31:16] = adder_tree_tier_6_p0_in[47:32] + adder_tree_tier_6_p0_in[63:48];
    adder_tree_tier_7_p0_in[47:32] = adder_tree_tier_6_p0_in[79:64] + adder_tree_tier_6_p0_in[95:80];
    adder_tree_tier_7_p0_in[63:48] = adder_tree_tier_6_p0_in[111:96];
    adder_tree_tier_8_p0_in[15:0] = adder_tree_tier_7_p0_in[15:0] + adder_tree_tier_7_p0_in[31:16];
    adder_tree_tier_8_p0_in[31:16] = adder_tree_tier_7_p0_in[47:32] + adder_tree_tier_7_p0_in[63:48];
    adder_tree_tier_9_p0_in[15:0] = adder_tree_tier_8_p0_in[15:0] + adder_tree_tier_8_p0_in[31:16];
    val_out_buffer[15:0] = adder_tree_tier_9_p0_in;
    adder_tree_tier_0_p1_in = tap_outputs[12831:6416];
    adder_tree_tier_1_p1_in[15:0] = adder_tree_tier_0_p1_in[15:0] + adder_tree_tier_0_p1_in[31:16];
    adder_tree_tier_1_p1_in[31:16] = adder_tree_tier_0_p1_in[47:32] + adder_tree_tier_0_p1_in[63:48];
    adder_tree_tier_1_p1_in[47:32] = adder_tree_tier_0_p1_in[79:64] + adder_tree_tier_0_p1_in[95:80];
    adder_tree_tier_1_p1_in[63:48] = adder_tree_tier_0_p1_in[111:96] + adder_tree_tier_0_p1_in[127:112];
    adder_tree_tier_1_p1_in[79:64] = adder_tree_tier_0_p1_in[143:128] + adder_tree_tier_0_p1_in[159:144];
    adder_tree_tier_1_p1_in[95:80] = adder_tree_tier_0_p1_in[175:160] + adder_tree_tier_0_p1_in[191:176];
    adder_tree_tier_1_p1_in[111:96] = adder_tree_tier_0_p1_in[207:192] + adder_tree_tier_0_p1_in[223:208];
    adder_tree_tier_1_p1_in[127:112] = adder_tree_tier_0_p1_in[239:224] + adder_tree_tier_0_p1_in[255:240];
    adder_tree_tier_1_p1_in[143:128] = adder_tree_tier_0_p1_in[271:256] + adder_tree_tier_0_p1_in[287:272];
    adder_tree_tier_1_p1_in[159:144] = adder_tree_tier_0_p1_in[303:288] + adder_tree_tier_0_p1_in[319:304];
    adder_tree_tier_1_p1_in[175:160] = adder_tree_tier_0_p1_in[335:320] + adder_tree_tier_0_p1_in[351:336];
    adder_tree_tier_1_p1_in[191:176] = adder_tree_tier_0_p1_in[367:352] + adder_tree_tier_0_p1_in[383:368];
    adder_tree_tier_1_p1_in[207:192] = adder_tree_tier_0_p1_in[399:384] + adder_tree_tier_0_p1_in[415:400];
    adder_tree_tier_1_p1_in[223:208] = adder_tree_tier_0_p1_in[431:416] + adder_tree_tier_0_p1_in[447:432];
    adder_tree_tier_1_p1_in[239:224] = adder_tree_tier_0_p1_in[463:448] + adder_tree_tier_0_p1_in[479:464];
    adder_tree_tier_1_p1_in[255:240] = adder_tree_tier_0_p1_in[495:480] + adder_tree_tier_0_p1_in[511:496];
    adder_tree_tier_1_p1_in[271:256] = adder_tree_tier_0_p1_in[527:512] + adder_tree_tier_0_p1_in[543:528];
    adder_tree_tier_1_p1_in[287:272] = adder_tree_tier_0_p1_in[559:544] + adder_tree_tier_0_p1_in[575:560];
    adder_tree_tier_1_p1_in[303:288] = adder_tree_tier_0_p1_in[591:576] + adder_tree_tier_0_p1_in[607:592];
    adder_tree_tier_1_p1_in[319:304] = adder_tree_tier_0_p1_in[623:608] + adder_tree_tier_0_p1_in[639:624];
    adder_tree_tier_1_p1_in[335:320] = adder_tree_tier_0_p1_in[655:640] + adder_tree_tier_0_p1_in[671:656];
    adder_tree_tier_1_p1_in[351:336] = adder_tree_tier_0_p1_in[687:672] + adder_tree_tier_0_p1_in[703:688];
    adder_tree_tier_1_p1_in[367:352] = adder_tree_tier_0_p1_in[719:704] + adder_tree_tier_0_p1_in[735:720];
    adder_tree_tier_1_p1_in[383:368] = adder_tree_tier_0_p1_in[751:736] + adder_tree_tier_0_p1_in[767:752];
    adder_tree_tier_1_p1_in[399:384] = adder_tree_tier_0_p1_in[783:768] + adder_tree_tier_0_p1_in[799:784];
    adder_tree_tier_1_p1_in[415:400] = adder_tree_tier_0_p1_in[815:800] + adder_tree_tier_0_p1_in[831:816];
    adder_tree_tier_1_p1_in[431:416] = adder_tree_tier_0_p1_in[847:832] + adder_tree_tier_0_p1_in[863:848];
    adder_tree_tier_1_p1_in[447:432] = adder_tree_tier_0_p1_in[879:864] + adder_tree_tier_0_p1_in[895:880];
    adder_tree_tier_1_p1_in[463:448] = adder_tree_tier_0_p1_in[911:896] + adder_tree_tier_0_p1_in[927:912];
    adder_tree_tier_1_p1_in[479:464] = adder_tree_tier_0_p1_in[943:928] + adder_tree_tier_0_p1_in[959:944];
    adder_tree_tier_1_p1_in[495:480] = adder_tree_tier_0_p1_in[975:960] + adder_tree_tier_0_p1_in[991:976];
    adder_tree_tier_1_p1_in[511:496] = adder_tree_tier_0_p1_in[1007:992] + adder_tree_tier_0_p1_in[1023:1008];
    adder_tree_tier_1_p1_in[527:512] = adder_tree_tier_0_p1_in[1039:1024] + adder_tree_tier_0_p1_in[1055:1040];
    adder_tree_tier_1_p1_in[543:528] = adder_tree_tier_0_p1_in[1071:1056] + adder_tree_tier_0_p1_in[1087:1072];
    adder_tree_tier_1_p1_in[559:544] = adder_tree_tier_0_p1_in[1103:1088] + adder_tree_tier_0_p1_in[1119:1104];
    adder_tree_tier_1_p1_in[575:560] = adder_tree_tier_0_p1_in[1135:1120] + adder_tree_tier_0_p1_in[1151:1136];
    adder_tree_tier_1_p1_in[591:576] = adder_tree_tier_0_p1_in[1167:1152] + adder_tree_tier_0_p1_in[1183:1168];
    adder_tree_tier_1_p1_in[607:592] = adder_tree_tier_0_p1_in[1199:1184] + adder_tree_tier_0_p1_in[1215:1200];
    adder_tree_tier_1_p1_in[623:608] = adder_tree_tier_0_p1_in[1231:1216] + adder_tree_tier_0_p1_in[1247:1232];
    adder_tree_tier_1_p1_in[639:624] = adder_tree_tier_0_p1_in[1263:1248] + adder_tree_tier_0_p1_in[1279:1264];
    adder_tree_tier_1_p1_in[655:640] = adder_tree_tier_0_p1_in[1295:1280] + adder_tree_tier_0_p1_in[1311:1296];
    adder_tree_tier_1_p1_in[671:656] = adder_tree_tier_0_p1_in[1327:1312] + adder_tree_tier_0_p1_in[1343:1328];
    adder_tree_tier_1_p1_in[687:672] = adder_tree_tier_0_p1_in[1359:1344] + adder_tree_tier_0_p1_in[1375:1360];
    adder_tree_tier_1_p1_in[703:688] = adder_tree_tier_0_p1_in[1391:1376] + adder_tree_tier_0_p1_in[1407:1392];
    adder_tree_tier_1_p1_in[719:704] = adder_tree_tier_0_p1_in[1423:1408] + adder_tree_tier_0_p1_in[1439:1424];
    adder_tree_tier_1_p1_in[735:720] = adder_tree_tier_0_p1_in[1455:1440] + adder_tree_tier_0_p1_in[1471:1456];
    adder_tree_tier_1_p1_in[751:736] = adder_tree_tier_0_p1_in[1487:1472] + adder_tree_tier_0_p1_in[1503:1488];
    adder_tree_tier_1_p1_in[767:752] = adder_tree_tier_0_p1_in[1519:1504] + adder_tree_tier_0_p1_in[1535:1520];
    adder_tree_tier_1_p1_in[783:768] = adder_tree_tier_0_p1_in[1551:1536] + adder_tree_tier_0_p1_in[1567:1552];
    adder_tree_tier_1_p1_in[799:784] = adder_tree_tier_0_p1_in[1583:1568] + adder_tree_tier_0_p1_in[1599:1584];
    adder_tree_tier_1_p1_in[815:800] = adder_tree_tier_0_p1_in[1615:1600] + adder_tree_tier_0_p1_in[1631:1616];
    adder_tree_tier_1_p1_in[831:816] = adder_tree_tier_0_p1_in[1647:1632] + adder_tree_tier_0_p1_in[1663:1648];
    adder_tree_tier_1_p1_in[847:832] = adder_tree_tier_0_p1_in[1679:1664] + adder_tree_tier_0_p1_in[1695:1680];
    adder_tree_tier_1_p1_in[863:848] = adder_tree_tier_0_p1_in[1711:1696] + adder_tree_tier_0_p1_in[1727:1712];
    adder_tree_tier_1_p1_in[879:864] = adder_tree_tier_0_p1_in[1743:1728] + adder_tree_tier_0_p1_in[1759:1744];
    adder_tree_tier_1_p1_in[895:880] = adder_tree_tier_0_p1_in[1775:1760] + adder_tree_tier_0_p1_in[1791:1776];
    adder_tree_tier_1_p1_in[911:896] = adder_tree_tier_0_p1_in[1807:1792] + adder_tree_tier_0_p1_in[1823:1808];
    adder_tree_tier_1_p1_in[927:912] = adder_tree_tier_0_p1_in[1839:1824] + adder_tree_tier_0_p1_in[1855:1840];
    adder_tree_tier_1_p1_in[943:928] = adder_tree_tier_0_p1_in[1871:1856] + adder_tree_tier_0_p1_in[1887:1872];
    adder_tree_tier_1_p1_in[959:944] = adder_tree_tier_0_p1_in[1903:1888] + adder_tree_tier_0_p1_in[1919:1904];
    adder_tree_tier_1_p1_in[975:960] = adder_tree_tier_0_p1_in[1935:1920] + adder_tree_tier_0_p1_in[1951:1936];
    adder_tree_tier_1_p1_in[991:976] = adder_tree_tier_0_p1_in[1967:1952] + adder_tree_tier_0_p1_in[1983:1968];
    adder_tree_tier_1_p1_in[1007:992] = adder_tree_tier_0_p1_in[1999:1984] + adder_tree_tier_0_p1_in[2015:2000];
    adder_tree_tier_1_p1_in[1023:1008] = adder_tree_tier_0_p1_in[2031:2016] + adder_tree_tier_0_p1_in[2047:2032];
    adder_tree_tier_1_p1_in[1039:1024] = adder_tree_tier_0_p1_in[2063:2048] + adder_tree_tier_0_p1_in[2079:2064];
    adder_tree_tier_1_p1_in[1055:1040] = adder_tree_tier_0_p1_in[2095:2080] + adder_tree_tier_0_p1_in[2111:2096];
    adder_tree_tier_1_p1_in[1071:1056] = adder_tree_tier_0_p1_in[2127:2112] + adder_tree_tier_0_p1_in[2143:2128];
    adder_tree_tier_1_p1_in[1087:1072] = adder_tree_tier_0_p1_in[2159:2144] + adder_tree_tier_0_p1_in[2175:2160];
    adder_tree_tier_1_p1_in[1103:1088] = adder_tree_tier_0_p1_in[2191:2176] + adder_tree_tier_0_p1_in[2207:2192];
    adder_tree_tier_1_p1_in[1119:1104] = adder_tree_tier_0_p1_in[2223:2208] + adder_tree_tier_0_p1_in[2239:2224];
    adder_tree_tier_1_p1_in[1135:1120] = adder_tree_tier_0_p1_in[2255:2240] + adder_tree_tier_0_p1_in[2271:2256];
    adder_tree_tier_1_p1_in[1151:1136] = adder_tree_tier_0_p1_in[2287:2272] + adder_tree_tier_0_p1_in[2303:2288];
    adder_tree_tier_1_p1_in[1167:1152] = adder_tree_tier_0_p1_in[2319:2304] + adder_tree_tier_0_p1_in[2335:2320];
    adder_tree_tier_1_p1_in[1183:1168] = adder_tree_tier_0_p1_in[2351:2336] + adder_tree_tier_0_p1_in[2367:2352];
    adder_tree_tier_1_p1_in[1199:1184] = adder_tree_tier_0_p1_in[2383:2368] + adder_tree_tier_0_p1_in[2399:2384];
    adder_tree_tier_1_p1_in[1215:1200] = adder_tree_tier_0_p1_in[2415:2400] + adder_tree_tier_0_p1_in[2431:2416];
    adder_tree_tier_1_p1_in[1231:1216] = adder_tree_tier_0_p1_in[2447:2432] + adder_tree_tier_0_p1_in[2463:2448];
    adder_tree_tier_1_p1_in[1247:1232] = adder_tree_tier_0_p1_in[2479:2464] + adder_tree_tier_0_p1_in[2495:2480];
    adder_tree_tier_1_p1_in[1263:1248] = adder_tree_tier_0_p1_in[2511:2496] + adder_tree_tier_0_p1_in[2527:2512];
    adder_tree_tier_1_p1_in[1279:1264] = adder_tree_tier_0_p1_in[2543:2528] + adder_tree_tier_0_p1_in[2559:2544];
    adder_tree_tier_1_p1_in[1295:1280] = adder_tree_tier_0_p1_in[2575:2560] + adder_tree_tier_0_p1_in[2591:2576];
    adder_tree_tier_1_p1_in[1311:1296] = adder_tree_tier_0_p1_in[2607:2592] + adder_tree_tier_0_p1_in[2623:2608];
    adder_tree_tier_1_p1_in[1327:1312] = adder_tree_tier_0_p1_in[2639:2624] + adder_tree_tier_0_p1_in[2655:2640];
    adder_tree_tier_1_p1_in[1343:1328] = adder_tree_tier_0_p1_in[2671:2656] + adder_tree_tier_0_p1_in[2687:2672];
    adder_tree_tier_1_p1_in[1359:1344] = adder_tree_tier_0_p1_in[2703:2688] + adder_tree_tier_0_p1_in[2719:2704];
    adder_tree_tier_1_p1_in[1375:1360] = adder_tree_tier_0_p1_in[2735:2720] + adder_tree_tier_0_p1_in[2751:2736];
    adder_tree_tier_1_p1_in[1391:1376] = adder_tree_tier_0_p1_in[2767:2752] + adder_tree_tier_0_p1_in[2783:2768];
    adder_tree_tier_1_p1_in[1407:1392] = adder_tree_tier_0_p1_in[2799:2784] + adder_tree_tier_0_p1_in[2815:2800];
    adder_tree_tier_1_p1_in[1423:1408] = adder_tree_tier_0_p1_in[2831:2816] + adder_tree_tier_0_p1_in[2847:2832];
    adder_tree_tier_1_p1_in[1439:1424] = adder_tree_tier_0_p1_in[2863:2848] + adder_tree_tier_0_p1_in[2879:2864];
    adder_tree_tier_1_p1_in[1455:1440] = adder_tree_tier_0_p1_in[2895:2880] + adder_tree_tier_0_p1_in[2911:2896];
    adder_tree_tier_1_p1_in[1471:1456] = adder_tree_tier_0_p1_in[2927:2912] + adder_tree_tier_0_p1_in[2943:2928];
    adder_tree_tier_1_p1_in[1487:1472] = adder_tree_tier_0_p1_in[2959:2944] + adder_tree_tier_0_p1_in[2975:2960];
    adder_tree_tier_1_p1_in[1503:1488] = adder_tree_tier_0_p1_in[2991:2976] + adder_tree_tier_0_p1_in[3007:2992];
    adder_tree_tier_1_p1_in[1519:1504] = adder_tree_tier_0_p1_in[3023:3008] + adder_tree_tier_0_p1_in[3039:3024];
    adder_tree_tier_1_p1_in[1535:1520] = adder_tree_tier_0_p1_in[3055:3040] + adder_tree_tier_0_p1_in[3071:3056];
    adder_tree_tier_1_p1_in[1551:1536] = adder_tree_tier_0_p1_in[3087:3072] + adder_tree_tier_0_p1_in[3103:3088];
    adder_tree_tier_1_p1_in[1567:1552] = adder_tree_tier_0_p1_in[3119:3104] + adder_tree_tier_0_p1_in[3135:3120];
    adder_tree_tier_1_p1_in[1583:1568] = adder_tree_tier_0_p1_in[3151:3136] + adder_tree_tier_0_p1_in[3167:3152];
    adder_tree_tier_1_p1_in[1599:1584] = adder_tree_tier_0_p1_in[3183:3168] + adder_tree_tier_0_p1_in[3199:3184];
    adder_tree_tier_1_p1_in[1615:1600] = adder_tree_tier_0_p1_in[3215:3200] + adder_tree_tier_0_p1_in[3231:3216];
    adder_tree_tier_1_p1_in[1631:1616] = adder_tree_tier_0_p1_in[3247:3232] + adder_tree_tier_0_p1_in[3263:3248];
    adder_tree_tier_1_p1_in[1647:1632] = adder_tree_tier_0_p1_in[3279:3264] + adder_tree_tier_0_p1_in[3295:3280];
    adder_tree_tier_1_p1_in[1663:1648] = adder_tree_tier_0_p1_in[3311:3296] + adder_tree_tier_0_p1_in[3327:3312];
    adder_tree_tier_1_p1_in[1679:1664] = adder_tree_tier_0_p1_in[3343:3328] + adder_tree_tier_0_p1_in[3359:3344];
    adder_tree_tier_1_p1_in[1695:1680] = adder_tree_tier_0_p1_in[3375:3360] + adder_tree_tier_0_p1_in[3391:3376];
    adder_tree_tier_1_p1_in[1711:1696] = adder_tree_tier_0_p1_in[3407:3392] + adder_tree_tier_0_p1_in[3423:3408];
    adder_tree_tier_1_p1_in[1727:1712] = adder_tree_tier_0_p1_in[3439:3424] + adder_tree_tier_0_p1_in[3455:3440];
    adder_tree_tier_1_p1_in[1743:1728] = adder_tree_tier_0_p1_in[3471:3456] + adder_tree_tier_0_p1_in[3487:3472];
    adder_tree_tier_1_p1_in[1759:1744] = adder_tree_tier_0_p1_in[3503:3488] + adder_tree_tier_0_p1_in[3519:3504];
    adder_tree_tier_1_p1_in[1775:1760] = adder_tree_tier_0_p1_in[3535:3520] + adder_tree_tier_0_p1_in[3551:3536];
    adder_tree_tier_1_p1_in[1791:1776] = adder_tree_tier_0_p1_in[3567:3552] + adder_tree_tier_0_p1_in[3583:3568];
    adder_tree_tier_1_p1_in[1807:1792] = adder_tree_tier_0_p1_in[3599:3584] + adder_tree_tier_0_p1_in[3615:3600];
    adder_tree_tier_1_p1_in[1823:1808] = adder_tree_tier_0_p1_in[3631:3616] + adder_tree_tier_0_p1_in[3647:3632];
    adder_tree_tier_1_p1_in[1839:1824] = adder_tree_tier_0_p1_in[3663:3648] + adder_tree_tier_0_p1_in[3679:3664];
    adder_tree_tier_1_p1_in[1855:1840] = adder_tree_tier_0_p1_in[3695:3680] + adder_tree_tier_0_p1_in[3711:3696];
    adder_tree_tier_1_p1_in[1871:1856] = adder_tree_tier_0_p1_in[3727:3712] + adder_tree_tier_0_p1_in[3743:3728];
    adder_tree_tier_1_p1_in[1887:1872] = adder_tree_tier_0_p1_in[3759:3744] + adder_tree_tier_0_p1_in[3775:3760];
    adder_tree_tier_1_p1_in[1903:1888] = adder_tree_tier_0_p1_in[3791:3776] + adder_tree_tier_0_p1_in[3807:3792];
    adder_tree_tier_1_p1_in[1919:1904] = adder_tree_tier_0_p1_in[3823:3808] + adder_tree_tier_0_p1_in[3839:3824];
    adder_tree_tier_1_p1_in[1935:1920] = adder_tree_tier_0_p1_in[3855:3840] + adder_tree_tier_0_p1_in[3871:3856];
    adder_tree_tier_1_p1_in[1951:1936] = adder_tree_tier_0_p1_in[3887:3872] + adder_tree_tier_0_p1_in[3903:3888];
    adder_tree_tier_1_p1_in[1967:1952] = adder_tree_tier_0_p1_in[3919:3904] + adder_tree_tier_0_p1_in[3935:3920];
    adder_tree_tier_1_p1_in[1983:1968] = adder_tree_tier_0_p1_in[3951:3936] + adder_tree_tier_0_p1_in[3967:3952];
    adder_tree_tier_1_p1_in[1999:1984] = adder_tree_tier_0_p1_in[3983:3968] + adder_tree_tier_0_p1_in[3999:3984];
    adder_tree_tier_1_p1_in[2015:2000] = adder_tree_tier_0_p1_in[4015:4000] + adder_tree_tier_0_p1_in[4031:4016];
    adder_tree_tier_1_p1_in[2031:2016] = adder_tree_tier_0_p1_in[4047:4032] + adder_tree_tier_0_p1_in[4063:4048];
    adder_tree_tier_1_p1_in[2047:2032] = adder_tree_tier_0_p1_in[4079:4064] + adder_tree_tier_0_p1_in[4095:4080];
    adder_tree_tier_1_p1_in[2063:2048] = adder_tree_tier_0_p1_in[4111:4096] + adder_tree_tier_0_p1_in[4127:4112];
    adder_tree_tier_1_p1_in[2079:2064] = adder_tree_tier_0_p1_in[4143:4128] + adder_tree_tier_0_p1_in[4159:4144];
    adder_tree_tier_1_p1_in[2095:2080] = adder_tree_tier_0_p1_in[4175:4160] + adder_tree_tier_0_p1_in[4191:4176];
    adder_tree_tier_1_p1_in[2111:2096] = adder_tree_tier_0_p1_in[4207:4192] + adder_tree_tier_0_p1_in[4223:4208];
    adder_tree_tier_1_p1_in[2127:2112] = adder_tree_tier_0_p1_in[4239:4224] + adder_tree_tier_0_p1_in[4255:4240];
    adder_tree_tier_1_p1_in[2143:2128] = adder_tree_tier_0_p1_in[4271:4256] + adder_tree_tier_0_p1_in[4287:4272];
    adder_tree_tier_1_p1_in[2159:2144] = adder_tree_tier_0_p1_in[4303:4288] + adder_tree_tier_0_p1_in[4319:4304];
    adder_tree_tier_1_p1_in[2175:2160] = adder_tree_tier_0_p1_in[4335:4320] + adder_tree_tier_0_p1_in[4351:4336];
    adder_tree_tier_1_p1_in[2191:2176] = adder_tree_tier_0_p1_in[4367:4352] + adder_tree_tier_0_p1_in[4383:4368];
    adder_tree_tier_1_p1_in[2207:2192] = adder_tree_tier_0_p1_in[4399:4384] + adder_tree_tier_0_p1_in[4415:4400];
    adder_tree_tier_1_p1_in[2223:2208] = adder_tree_tier_0_p1_in[4431:4416] + adder_tree_tier_0_p1_in[4447:4432];
    adder_tree_tier_1_p1_in[2239:2224] = adder_tree_tier_0_p1_in[4463:4448] + adder_tree_tier_0_p1_in[4479:4464];
    adder_tree_tier_1_p1_in[2255:2240] = adder_tree_tier_0_p1_in[4495:4480] + adder_tree_tier_0_p1_in[4511:4496];
    adder_tree_tier_1_p1_in[2271:2256] = adder_tree_tier_0_p1_in[4527:4512] + adder_tree_tier_0_p1_in[4543:4528];
    adder_tree_tier_1_p1_in[2287:2272] = adder_tree_tier_0_p1_in[4559:4544] + adder_tree_tier_0_p1_in[4575:4560];
    adder_tree_tier_1_p1_in[2303:2288] = adder_tree_tier_0_p1_in[4591:4576] + adder_tree_tier_0_p1_in[4607:4592];
    adder_tree_tier_1_p1_in[2319:2304] = adder_tree_tier_0_p1_in[4623:4608] + adder_tree_tier_0_p1_in[4639:4624];
    adder_tree_tier_1_p1_in[2335:2320] = adder_tree_tier_0_p1_in[4655:4640] + adder_tree_tier_0_p1_in[4671:4656];
    adder_tree_tier_1_p1_in[2351:2336] = adder_tree_tier_0_p1_in[4687:4672] + adder_tree_tier_0_p1_in[4703:4688];
    adder_tree_tier_1_p1_in[2367:2352] = adder_tree_tier_0_p1_in[4719:4704] + adder_tree_tier_0_p1_in[4735:4720];
    adder_tree_tier_1_p1_in[2383:2368] = adder_tree_tier_0_p1_in[4751:4736] + adder_tree_tier_0_p1_in[4767:4752];
    adder_tree_tier_1_p1_in[2399:2384] = adder_tree_tier_0_p1_in[4783:4768] + adder_tree_tier_0_p1_in[4799:4784];
    adder_tree_tier_1_p1_in[2415:2400] = adder_tree_tier_0_p1_in[4815:4800] + adder_tree_tier_0_p1_in[4831:4816];
    adder_tree_tier_1_p1_in[2431:2416] = adder_tree_tier_0_p1_in[4847:4832] + adder_tree_tier_0_p1_in[4863:4848];
    adder_tree_tier_1_p1_in[2447:2432] = adder_tree_tier_0_p1_in[4879:4864] + adder_tree_tier_0_p1_in[4895:4880];
    adder_tree_tier_1_p1_in[2463:2448] = adder_tree_tier_0_p1_in[4911:4896] + adder_tree_tier_0_p1_in[4927:4912];
    adder_tree_tier_1_p1_in[2479:2464] = adder_tree_tier_0_p1_in[4943:4928] + adder_tree_tier_0_p1_in[4959:4944];
    adder_tree_tier_1_p1_in[2495:2480] = adder_tree_tier_0_p1_in[4975:4960] + adder_tree_tier_0_p1_in[4991:4976];
    adder_tree_tier_1_p1_in[2511:2496] = adder_tree_tier_0_p1_in[5007:4992] + adder_tree_tier_0_p1_in[5023:5008];
    adder_tree_tier_1_p1_in[2527:2512] = adder_tree_tier_0_p1_in[5039:5024] + adder_tree_tier_0_p1_in[5055:5040];
    adder_tree_tier_1_p1_in[2543:2528] = adder_tree_tier_0_p1_in[5071:5056] + adder_tree_tier_0_p1_in[5087:5072];
    adder_tree_tier_1_p1_in[2559:2544] = adder_tree_tier_0_p1_in[5103:5088] + adder_tree_tier_0_p1_in[5119:5104];
    adder_tree_tier_1_p1_in[2575:2560] = adder_tree_tier_0_p1_in[5135:5120] + adder_tree_tier_0_p1_in[5151:5136];
    adder_tree_tier_1_p1_in[2591:2576] = adder_tree_tier_0_p1_in[5167:5152] + adder_tree_tier_0_p1_in[5183:5168];
    adder_tree_tier_1_p1_in[2607:2592] = adder_tree_tier_0_p1_in[5199:5184] + adder_tree_tier_0_p1_in[5215:5200];
    adder_tree_tier_1_p1_in[2623:2608] = adder_tree_tier_0_p1_in[5231:5216] + adder_tree_tier_0_p1_in[5247:5232];
    adder_tree_tier_1_p1_in[2639:2624] = adder_tree_tier_0_p1_in[5263:5248] + adder_tree_tier_0_p1_in[5279:5264];
    adder_tree_tier_1_p1_in[2655:2640] = adder_tree_tier_0_p1_in[5295:5280] + adder_tree_tier_0_p1_in[5311:5296];
    adder_tree_tier_1_p1_in[2671:2656] = adder_tree_tier_0_p1_in[5327:5312] + adder_tree_tier_0_p1_in[5343:5328];
    adder_tree_tier_1_p1_in[2687:2672] = adder_tree_tier_0_p1_in[5359:5344] + adder_tree_tier_0_p1_in[5375:5360];
    adder_tree_tier_1_p1_in[2703:2688] = adder_tree_tier_0_p1_in[5391:5376] + adder_tree_tier_0_p1_in[5407:5392];
    adder_tree_tier_1_p1_in[2719:2704] = adder_tree_tier_0_p1_in[5423:5408] + adder_tree_tier_0_p1_in[5439:5424];
    adder_tree_tier_1_p1_in[2735:2720] = adder_tree_tier_0_p1_in[5455:5440] + adder_tree_tier_0_p1_in[5471:5456];
    adder_tree_tier_1_p1_in[2751:2736] = adder_tree_tier_0_p1_in[5487:5472] + adder_tree_tier_0_p1_in[5503:5488];
    adder_tree_tier_1_p1_in[2767:2752] = adder_tree_tier_0_p1_in[5519:5504] + adder_tree_tier_0_p1_in[5535:5520];
    adder_tree_tier_1_p1_in[2783:2768] = adder_tree_tier_0_p1_in[5551:5536] + adder_tree_tier_0_p1_in[5567:5552];
    adder_tree_tier_1_p1_in[2799:2784] = adder_tree_tier_0_p1_in[5583:5568] + adder_tree_tier_0_p1_in[5599:5584];
    adder_tree_tier_1_p1_in[2815:2800] = adder_tree_tier_0_p1_in[5615:5600] + adder_tree_tier_0_p1_in[5631:5616];
    adder_tree_tier_1_p1_in[2831:2816] = adder_tree_tier_0_p1_in[5647:5632] + adder_tree_tier_0_p1_in[5663:5648];
    adder_tree_tier_1_p1_in[2847:2832] = adder_tree_tier_0_p1_in[5679:5664] + adder_tree_tier_0_p1_in[5695:5680];
    adder_tree_tier_1_p1_in[2863:2848] = adder_tree_tier_0_p1_in[5711:5696] + adder_tree_tier_0_p1_in[5727:5712];
    adder_tree_tier_1_p1_in[2879:2864] = adder_tree_tier_0_p1_in[5743:5728] + adder_tree_tier_0_p1_in[5759:5744];
    adder_tree_tier_1_p1_in[2895:2880] = adder_tree_tier_0_p1_in[5775:5760] + adder_tree_tier_0_p1_in[5791:5776];
    adder_tree_tier_1_p1_in[2911:2896] = adder_tree_tier_0_p1_in[5807:5792] + adder_tree_tier_0_p1_in[5823:5808];
    adder_tree_tier_1_p1_in[2927:2912] = adder_tree_tier_0_p1_in[5839:5824] + adder_tree_tier_0_p1_in[5855:5840];
    adder_tree_tier_1_p1_in[2943:2928] = adder_tree_tier_0_p1_in[5871:5856] + adder_tree_tier_0_p1_in[5887:5872];
    adder_tree_tier_1_p1_in[2959:2944] = adder_tree_tier_0_p1_in[5903:5888] + adder_tree_tier_0_p1_in[5919:5904];
    adder_tree_tier_1_p1_in[2975:2960] = adder_tree_tier_0_p1_in[5935:5920] + adder_tree_tier_0_p1_in[5951:5936];
    adder_tree_tier_1_p1_in[2991:2976] = adder_tree_tier_0_p1_in[5967:5952] + adder_tree_tier_0_p1_in[5983:5968];
    adder_tree_tier_1_p1_in[3007:2992] = adder_tree_tier_0_p1_in[5999:5984] + adder_tree_tier_0_p1_in[6015:6000];
    adder_tree_tier_1_p1_in[3023:3008] = adder_tree_tier_0_p1_in[6031:6016] + adder_tree_tier_0_p1_in[6047:6032];
    adder_tree_tier_1_p1_in[3039:3024] = adder_tree_tier_0_p1_in[6063:6048] + adder_tree_tier_0_p1_in[6079:6064];
    adder_tree_tier_1_p1_in[3055:3040] = adder_tree_tier_0_p1_in[6095:6080] + adder_tree_tier_0_p1_in[6111:6096];
    adder_tree_tier_1_p1_in[3071:3056] = adder_tree_tier_0_p1_in[6127:6112] + adder_tree_tier_0_p1_in[6143:6128];
    adder_tree_tier_1_p1_in[3087:3072] = adder_tree_tier_0_p1_in[6159:6144] + adder_tree_tier_0_p1_in[6175:6160];
    adder_tree_tier_1_p1_in[3103:3088] = adder_tree_tier_0_p1_in[6191:6176] + adder_tree_tier_0_p1_in[6207:6192];
    adder_tree_tier_1_p1_in[3119:3104] = adder_tree_tier_0_p1_in[6223:6208] + adder_tree_tier_0_p1_in[6239:6224];
    adder_tree_tier_1_p1_in[3135:3120] = adder_tree_tier_0_p1_in[6255:6240] + adder_tree_tier_0_p1_in[6271:6256];
    adder_tree_tier_1_p1_in[3151:3136] = adder_tree_tier_0_p1_in[6287:6272] + adder_tree_tier_0_p1_in[6303:6288];
    adder_tree_tier_1_p1_in[3167:3152] = adder_tree_tier_0_p1_in[6319:6304] + adder_tree_tier_0_p1_in[6335:6320];
    adder_tree_tier_1_p1_in[3183:3168] = adder_tree_tier_0_p1_in[6351:6336] + adder_tree_tier_0_p1_in[6367:6352];
    adder_tree_tier_1_p1_in[3199:3184] = adder_tree_tier_0_p1_in[6383:6368] + adder_tree_tier_0_p1_in[6399:6384];
    adder_tree_tier_1_p1_in[3215:3200] = adder_tree_tier_0_p1_in[6415:6400];
    adder_tree_tier_2_p1_in[15:0] = adder_tree_tier_1_p1_in[15:0] + adder_tree_tier_1_p1_in[31:16];
    adder_tree_tier_2_p1_in[31:16] = adder_tree_tier_1_p1_in[47:32] + adder_tree_tier_1_p1_in[63:48];
    adder_tree_tier_2_p1_in[47:32] = adder_tree_tier_1_p1_in[79:64] + adder_tree_tier_1_p1_in[95:80];
    adder_tree_tier_2_p1_in[63:48] = adder_tree_tier_1_p1_in[111:96] + adder_tree_tier_1_p1_in[127:112];
    adder_tree_tier_2_p1_in[79:64] = adder_tree_tier_1_p1_in[143:128] + adder_tree_tier_1_p1_in[159:144];
    adder_tree_tier_2_p1_in[95:80] = adder_tree_tier_1_p1_in[175:160] + adder_tree_tier_1_p1_in[191:176];
    adder_tree_tier_2_p1_in[111:96] = adder_tree_tier_1_p1_in[207:192] + adder_tree_tier_1_p1_in[223:208];
    adder_tree_tier_2_p1_in[127:112] = adder_tree_tier_1_p1_in[239:224] + adder_tree_tier_1_p1_in[255:240];
    adder_tree_tier_2_p1_in[143:128] = adder_tree_tier_1_p1_in[271:256] + adder_tree_tier_1_p1_in[287:272];
    adder_tree_tier_2_p1_in[159:144] = adder_tree_tier_1_p1_in[303:288] + adder_tree_tier_1_p1_in[319:304];
    adder_tree_tier_2_p1_in[175:160] = adder_tree_tier_1_p1_in[335:320] + adder_tree_tier_1_p1_in[351:336];
    adder_tree_tier_2_p1_in[191:176] = adder_tree_tier_1_p1_in[367:352] + adder_tree_tier_1_p1_in[383:368];
    adder_tree_tier_2_p1_in[207:192] = adder_tree_tier_1_p1_in[399:384] + adder_tree_tier_1_p1_in[415:400];
    adder_tree_tier_2_p1_in[223:208] = adder_tree_tier_1_p1_in[431:416] + adder_tree_tier_1_p1_in[447:432];
    adder_tree_tier_2_p1_in[239:224] = adder_tree_tier_1_p1_in[463:448] + adder_tree_tier_1_p1_in[479:464];
    adder_tree_tier_2_p1_in[255:240] = adder_tree_tier_1_p1_in[495:480] + adder_tree_tier_1_p1_in[511:496];
    adder_tree_tier_2_p1_in[271:256] = adder_tree_tier_1_p1_in[527:512] + adder_tree_tier_1_p1_in[543:528];
    adder_tree_tier_2_p1_in[287:272] = adder_tree_tier_1_p1_in[559:544] + adder_tree_tier_1_p1_in[575:560];
    adder_tree_tier_2_p1_in[303:288] = adder_tree_tier_1_p1_in[591:576] + adder_tree_tier_1_p1_in[607:592];
    adder_tree_tier_2_p1_in[319:304] = adder_tree_tier_1_p1_in[623:608] + adder_tree_tier_1_p1_in[639:624];
    adder_tree_tier_2_p1_in[335:320] = adder_tree_tier_1_p1_in[655:640] + adder_tree_tier_1_p1_in[671:656];
    adder_tree_tier_2_p1_in[351:336] = adder_tree_tier_1_p1_in[687:672] + adder_tree_tier_1_p1_in[703:688];
    adder_tree_tier_2_p1_in[367:352] = adder_tree_tier_1_p1_in[719:704] + adder_tree_tier_1_p1_in[735:720];
    adder_tree_tier_2_p1_in[383:368] = adder_tree_tier_1_p1_in[751:736] + adder_tree_tier_1_p1_in[767:752];
    adder_tree_tier_2_p1_in[399:384] = adder_tree_tier_1_p1_in[783:768] + adder_tree_tier_1_p1_in[799:784];
    adder_tree_tier_2_p1_in[415:400] = adder_tree_tier_1_p1_in[815:800] + adder_tree_tier_1_p1_in[831:816];
    adder_tree_tier_2_p1_in[431:416] = adder_tree_tier_1_p1_in[847:832] + adder_tree_tier_1_p1_in[863:848];
    adder_tree_tier_2_p1_in[447:432] = adder_tree_tier_1_p1_in[879:864] + adder_tree_tier_1_p1_in[895:880];
    adder_tree_tier_2_p1_in[463:448] = adder_tree_tier_1_p1_in[911:896] + adder_tree_tier_1_p1_in[927:912];
    adder_tree_tier_2_p1_in[479:464] = adder_tree_tier_1_p1_in[943:928] + adder_tree_tier_1_p1_in[959:944];
    adder_tree_tier_2_p1_in[495:480] = adder_tree_tier_1_p1_in[975:960] + adder_tree_tier_1_p1_in[991:976];
    adder_tree_tier_2_p1_in[511:496] = adder_tree_tier_1_p1_in[1007:992] + adder_tree_tier_1_p1_in[1023:1008];
    adder_tree_tier_2_p1_in[527:512] = adder_tree_tier_1_p1_in[1039:1024] + adder_tree_tier_1_p1_in[1055:1040];
    adder_tree_tier_2_p1_in[543:528] = adder_tree_tier_1_p1_in[1071:1056] + adder_tree_tier_1_p1_in[1087:1072];
    adder_tree_tier_2_p1_in[559:544] = adder_tree_tier_1_p1_in[1103:1088] + adder_tree_tier_1_p1_in[1119:1104];
    adder_tree_tier_2_p1_in[575:560] = adder_tree_tier_1_p1_in[1135:1120] + adder_tree_tier_1_p1_in[1151:1136];
    adder_tree_tier_2_p1_in[591:576] = adder_tree_tier_1_p1_in[1167:1152] + adder_tree_tier_1_p1_in[1183:1168];
    adder_tree_tier_2_p1_in[607:592] = adder_tree_tier_1_p1_in[1199:1184] + adder_tree_tier_1_p1_in[1215:1200];
    adder_tree_tier_2_p1_in[623:608] = adder_tree_tier_1_p1_in[1231:1216] + adder_tree_tier_1_p1_in[1247:1232];
    adder_tree_tier_2_p1_in[639:624] = adder_tree_tier_1_p1_in[1263:1248] + adder_tree_tier_1_p1_in[1279:1264];
    adder_tree_tier_2_p1_in[655:640] = adder_tree_tier_1_p1_in[1295:1280] + adder_tree_tier_1_p1_in[1311:1296];
    adder_tree_tier_2_p1_in[671:656] = adder_tree_tier_1_p1_in[1327:1312] + adder_tree_tier_1_p1_in[1343:1328];
    adder_tree_tier_2_p1_in[687:672] = adder_tree_tier_1_p1_in[1359:1344] + adder_tree_tier_1_p1_in[1375:1360];
    adder_tree_tier_2_p1_in[703:688] = adder_tree_tier_1_p1_in[1391:1376] + adder_tree_tier_1_p1_in[1407:1392];
    adder_tree_tier_2_p1_in[719:704] = adder_tree_tier_1_p1_in[1423:1408] + adder_tree_tier_1_p1_in[1439:1424];
    adder_tree_tier_2_p1_in[735:720] = adder_tree_tier_1_p1_in[1455:1440] + adder_tree_tier_1_p1_in[1471:1456];
    adder_tree_tier_2_p1_in[751:736] = adder_tree_tier_1_p1_in[1487:1472] + adder_tree_tier_1_p1_in[1503:1488];
    adder_tree_tier_2_p1_in[767:752] = adder_tree_tier_1_p1_in[1519:1504] + adder_tree_tier_1_p1_in[1535:1520];
    adder_tree_tier_2_p1_in[783:768] = adder_tree_tier_1_p1_in[1551:1536] + adder_tree_tier_1_p1_in[1567:1552];
    adder_tree_tier_2_p1_in[799:784] = adder_tree_tier_1_p1_in[1583:1568] + adder_tree_tier_1_p1_in[1599:1584];
    adder_tree_tier_2_p1_in[815:800] = adder_tree_tier_1_p1_in[1615:1600] + adder_tree_tier_1_p1_in[1631:1616];
    adder_tree_tier_2_p1_in[831:816] = adder_tree_tier_1_p1_in[1647:1632] + adder_tree_tier_1_p1_in[1663:1648];
    adder_tree_tier_2_p1_in[847:832] = adder_tree_tier_1_p1_in[1679:1664] + adder_tree_tier_1_p1_in[1695:1680];
    adder_tree_tier_2_p1_in[863:848] = adder_tree_tier_1_p1_in[1711:1696] + adder_tree_tier_1_p1_in[1727:1712];
    adder_tree_tier_2_p1_in[879:864] = adder_tree_tier_1_p1_in[1743:1728] + adder_tree_tier_1_p1_in[1759:1744];
    adder_tree_tier_2_p1_in[895:880] = adder_tree_tier_1_p1_in[1775:1760] + adder_tree_tier_1_p1_in[1791:1776];
    adder_tree_tier_2_p1_in[911:896] = adder_tree_tier_1_p1_in[1807:1792] + adder_tree_tier_1_p1_in[1823:1808];
    adder_tree_tier_2_p1_in[927:912] = adder_tree_tier_1_p1_in[1839:1824] + adder_tree_tier_1_p1_in[1855:1840];
    adder_tree_tier_2_p1_in[943:928] = adder_tree_tier_1_p1_in[1871:1856] + adder_tree_tier_1_p1_in[1887:1872];
    adder_tree_tier_2_p1_in[959:944] = adder_tree_tier_1_p1_in[1903:1888] + adder_tree_tier_1_p1_in[1919:1904];
    adder_tree_tier_2_p1_in[975:960] = adder_tree_tier_1_p1_in[1935:1920] + adder_tree_tier_1_p1_in[1951:1936];
    adder_tree_tier_2_p1_in[991:976] = adder_tree_tier_1_p1_in[1967:1952] + adder_tree_tier_1_p1_in[1983:1968];
    adder_tree_tier_2_p1_in[1007:992] = adder_tree_tier_1_p1_in[1999:1984] + adder_tree_tier_1_p1_in[2015:2000];
    adder_tree_tier_2_p1_in[1023:1008] = adder_tree_tier_1_p1_in[2031:2016] + adder_tree_tier_1_p1_in[2047:2032];
    adder_tree_tier_2_p1_in[1039:1024] = adder_tree_tier_1_p1_in[2063:2048] + adder_tree_tier_1_p1_in[2079:2064];
    adder_tree_tier_2_p1_in[1055:1040] = adder_tree_tier_1_p1_in[2095:2080] + adder_tree_tier_1_p1_in[2111:2096];
    adder_tree_tier_2_p1_in[1071:1056] = adder_tree_tier_1_p1_in[2127:2112] + adder_tree_tier_1_p1_in[2143:2128];
    adder_tree_tier_2_p1_in[1087:1072] = adder_tree_tier_1_p1_in[2159:2144] + adder_tree_tier_1_p1_in[2175:2160];
    adder_tree_tier_2_p1_in[1103:1088] = adder_tree_tier_1_p1_in[2191:2176] + adder_tree_tier_1_p1_in[2207:2192];
    adder_tree_tier_2_p1_in[1119:1104] = adder_tree_tier_1_p1_in[2223:2208] + adder_tree_tier_1_p1_in[2239:2224];
    adder_tree_tier_2_p1_in[1135:1120] = adder_tree_tier_1_p1_in[2255:2240] + adder_tree_tier_1_p1_in[2271:2256];
    adder_tree_tier_2_p1_in[1151:1136] = adder_tree_tier_1_p1_in[2287:2272] + adder_tree_tier_1_p1_in[2303:2288];
    adder_tree_tier_2_p1_in[1167:1152] = adder_tree_tier_1_p1_in[2319:2304] + adder_tree_tier_1_p1_in[2335:2320];
    adder_tree_tier_2_p1_in[1183:1168] = adder_tree_tier_1_p1_in[2351:2336] + adder_tree_tier_1_p1_in[2367:2352];
    adder_tree_tier_2_p1_in[1199:1184] = adder_tree_tier_1_p1_in[2383:2368] + adder_tree_tier_1_p1_in[2399:2384];
    adder_tree_tier_2_p1_in[1215:1200] = adder_tree_tier_1_p1_in[2415:2400] + adder_tree_tier_1_p1_in[2431:2416];
    adder_tree_tier_2_p1_in[1231:1216] = adder_tree_tier_1_p1_in[2447:2432] + adder_tree_tier_1_p1_in[2463:2448];
    adder_tree_tier_2_p1_in[1247:1232] = adder_tree_tier_1_p1_in[2479:2464] + adder_tree_tier_1_p1_in[2495:2480];
    adder_tree_tier_2_p1_in[1263:1248] = adder_tree_tier_1_p1_in[2511:2496] + adder_tree_tier_1_p1_in[2527:2512];
    adder_tree_tier_2_p1_in[1279:1264] = adder_tree_tier_1_p1_in[2543:2528] + adder_tree_tier_1_p1_in[2559:2544];
    adder_tree_tier_2_p1_in[1295:1280] = adder_tree_tier_1_p1_in[2575:2560] + adder_tree_tier_1_p1_in[2591:2576];
    adder_tree_tier_2_p1_in[1311:1296] = adder_tree_tier_1_p1_in[2607:2592] + adder_tree_tier_1_p1_in[2623:2608];
    adder_tree_tier_2_p1_in[1327:1312] = adder_tree_tier_1_p1_in[2639:2624] + adder_tree_tier_1_p1_in[2655:2640];
    adder_tree_tier_2_p1_in[1343:1328] = adder_tree_tier_1_p1_in[2671:2656] + adder_tree_tier_1_p1_in[2687:2672];
    adder_tree_tier_2_p1_in[1359:1344] = adder_tree_tier_1_p1_in[2703:2688] + adder_tree_tier_1_p1_in[2719:2704];
    adder_tree_tier_2_p1_in[1375:1360] = adder_tree_tier_1_p1_in[2735:2720] + adder_tree_tier_1_p1_in[2751:2736];
    adder_tree_tier_2_p1_in[1391:1376] = adder_tree_tier_1_p1_in[2767:2752] + adder_tree_tier_1_p1_in[2783:2768];
    adder_tree_tier_2_p1_in[1407:1392] = adder_tree_tier_1_p1_in[2799:2784] + adder_tree_tier_1_p1_in[2815:2800];
    adder_tree_tier_2_p1_in[1423:1408] = adder_tree_tier_1_p1_in[2831:2816] + adder_tree_tier_1_p1_in[2847:2832];
    adder_tree_tier_2_p1_in[1439:1424] = adder_tree_tier_1_p1_in[2863:2848] + adder_tree_tier_1_p1_in[2879:2864];
    adder_tree_tier_2_p1_in[1455:1440] = adder_tree_tier_1_p1_in[2895:2880] + adder_tree_tier_1_p1_in[2911:2896];
    adder_tree_tier_2_p1_in[1471:1456] = adder_tree_tier_1_p1_in[2927:2912] + adder_tree_tier_1_p1_in[2943:2928];
    adder_tree_tier_2_p1_in[1487:1472] = adder_tree_tier_1_p1_in[2959:2944] + adder_tree_tier_1_p1_in[2975:2960];
    adder_tree_tier_2_p1_in[1503:1488] = adder_tree_tier_1_p1_in[2991:2976] + adder_tree_tier_1_p1_in[3007:2992];
    adder_tree_tier_2_p1_in[1519:1504] = adder_tree_tier_1_p1_in[3023:3008] + adder_tree_tier_1_p1_in[3039:3024];
    adder_tree_tier_2_p1_in[1535:1520] = adder_tree_tier_1_p1_in[3055:3040] + adder_tree_tier_1_p1_in[3071:3056];
    adder_tree_tier_2_p1_in[1551:1536] = adder_tree_tier_1_p1_in[3087:3072] + adder_tree_tier_1_p1_in[3103:3088];
    adder_tree_tier_2_p1_in[1567:1552] = adder_tree_tier_1_p1_in[3119:3104] + adder_tree_tier_1_p1_in[3135:3120];
    adder_tree_tier_2_p1_in[1583:1568] = adder_tree_tier_1_p1_in[3151:3136] + adder_tree_tier_1_p1_in[3167:3152];
    adder_tree_tier_2_p1_in[1599:1584] = adder_tree_tier_1_p1_in[3183:3168] + adder_tree_tier_1_p1_in[3199:3184];
    adder_tree_tier_2_p1_in[1615:1600] = adder_tree_tier_1_p1_in[3215:3200];
    adder_tree_tier_3_p1_in[15:0] = adder_tree_tier_2_p1_in[15:0] + adder_tree_tier_2_p1_in[31:16];
    adder_tree_tier_3_p1_in[31:16] = adder_tree_tier_2_p1_in[47:32] + adder_tree_tier_2_p1_in[63:48];
    adder_tree_tier_3_p1_in[47:32] = adder_tree_tier_2_p1_in[79:64] + adder_tree_tier_2_p1_in[95:80];
    adder_tree_tier_3_p1_in[63:48] = adder_tree_tier_2_p1_in[111:96] + adder_tree_tier_2_p1_in[127:112];
    adder_tree_tier_3_p1_in[79:64] = adder_tree_tier_2_p1_in[143:128] + adder_tree_tier_2_p1_in[159:144];
    adder_tree_tier_3_p1_in[95:80] = adder_tree_tier_2_p1_in[175:160] + adder_tree_tier_2_p1_in[191:176];
    adder_tree_tier_3_p1_in[111:96] = adder_tree_tier_2_p1_in[207:192] + adder_tree_tier_2_p1_in[223:208];
    adder_tree_tier_3_p1_in[127:112] = adder_tree_tier_2_p1_in[239:224] + adder_tree_tier_2_p1_in[255:240];
    adder_tree_tier_3_p1_in[143:128] = adder_tree_tier_2_p1_in[271:256] + adder_tree_tier_2_p1_in[287:272];
    adder_tree_tier_3_p1_in[159:144] = adder_tree_tier_2_p1_in[303:288] + adder_tree_tier_2_p1_in[319:304];
    adder_tree_tier_3_p1_in[175:160] = adder_tree_tier_2_p1_in[335:320] + adder_tree_tier_2_p1_in[351:336];
    adder_tree_tier_3_p1_in[191:176] = adder_tree_tier_2_p1_in[367:352] + adder_tree_tier_2_p1_in[383:368];
    adder_tree_tier_3_p1_in[207:192] = adder_tree_tier_2_p1_in[399:384] + adder_tree_tier_2_p1_in[415:400];
    adder_tree_tier_3_p1_in[223:208] = adder_tree_tier_2_p1_in[431:416] + adder_tree_tier_2_p1_in[447:432];
    adder_tree_tier_3_p1_in[239:224] = adder_tree_tier_2_p1_in[463:448] + adder_tree_tier_2_p1_in[479:464];
    adder_tree_tier_3_p1_in[255:240] = adder_tree_tier_2_p1_in[495:480] + adder_tree_tier_2_p1_in[511:496];
    adder_tree_tier_3_p1_in[271:256] = adder_tree_tier_2_p1_in[527:512] + adder_tree_tier_2_p1_in[543:528];
    adder_tree_tier_3_p1_in[287:272] = adder_tree_tier_2_p1_in[559:544] + adder_tree_tier_2_p1_in[575:560];
    adder_tree_tier_3_p1_in[303:288] = adder_tree_tier_2_p1_in[591:576] + adder_tree_tier_2_p1_in[607:592];
    adder_tree_tier_3_p1_in[319:304] = adder_tree_tier_2_p1_in[623:608] + adder_tree_tier_2_p1_in[639:624];
    adder_tree_tier_3_p1_in[335:320] = adder_tree_tier_2_p1_in[655:640] + adder_tree_tier_2_p1_in[671:656];
    adder_tree_tier_3_p1_in[351:336] = adder_tree_tier_2_p1_in[687:672] + adder_tree_tier_2_p1_in[703:688];
    adder_tree_tier_3_p1_in[367:352] = adder_tree_tier_2_p1_in[719:704] + adder_tree_tier_2_p1_in[735:720];
    adder_tree_tier_3_p1_in[383:368] = adder_tree_tier_2_p1_in[751:736] + adder_tree_tier_2_p1_in[767:752];
    adder_tree_tier_3_p1_in[399:384] = adder_tree_tier_2_p1_in[783:768] + adder_tree_tier_2_p1_in[799:784];
    adder_tree_tier_3_p1_in[415:400] = adder_tree_tier_2_p1_in[815:800] + adder_tree_tier_2_p1_in[831:816];
    adder_tree_tier_3_p1_in[431:416] = adder_tree_tier_2_p1_in[847:832] + adder_tree_tier_2_p1_in[863:848];
    adder_tree_tier_3_p1_in[447:432] = adder_tree_tier_2_p1_in[879:864] + adder_tree_tier_2_p1_in[895:880];
    adder_tree_tier_3_p1_in[463:448] = adder_tree_tier_2_p1_in[911:896] + adder_tree_tier_2_p1_in[927:912];
    adder_tree_tier_3_p1_in[479:464] = adder_tree_tier_2_p1_in[943:928] + adder_tree_tier_2_p1_in[959:944];
    adder_tree_tier_3_p1_in[495:480] = adder_tree_tier_2_p1_in[975:960] + adder_tree_tier_2_p1_in[991:976];
    adder_tree_tier_3_p1_in[511:496] = adder_tree_tier_2_p1_in[1007:992] + adder_tree_tier_2_p1_in[1023:1008];
    adder_tree_tier_3_p1_in[527:512] = adder_tree_tier_2_p1_in[1039:1024] + adder_tree_tier_2_p1_in[1055:1040];
    adder_tree_tier_3_p1_in[543:528] = adder_tree_tier_2_p1_in[1071:1056] + adder_tree_tier_2_p1_in[1087:1072];
    adder_tree_tier_3_p1_in[559:544] = adder_tree_tier_2_p1_in[1103:1088] + adder_tree_tier_2_p1_in[1119:1104];
    adder_tree_tier_3_p1_in[575:560] = adder_tree_tier_2_p1_in[1135:1120] + adder_tree_tier_2_p1_in[1151:1136];
    adder_tree_tier_3_p1_in[591:576] = adder_tree_tier_2_p1_in[1167:1152] + adder_tree_tier_2_p1_in[1183:1168];
    adder_tree_tier_3_p1_in[607:592] = adder_tree_tier_2_p1_in[1199:1184] + adder_tree_tier_2_p1_in[1215:1200];
    adder_tree_tier_3_p1_in[623:608] = adder_tree_tier_2_p1_in[1231:1216] + adder_tree_tier_2_p1_in[1247:1232];
    adder_tree_tier_3_p1_in[639:624] = adder_tree_tier_2_p1_in[1263:1248] + adder_tree_tier_2_p1_in[1279:1264];
    adder_tree_tier_3_p1_in[655:640] = adder_tree_tier_2_p1_in[1295:1280] + adder_tree_tier_2_p1_in[1311:1296];
    adder_tree_tier_3_p1_in[671:656] = adder_tree_tier_2_p1_in[1327:1312] + adder_tree_tier_2_p1_in[1343:1328];
    adder_tree_tier_3_p1_in[687:672] = adder_tree_tier_2_p1_in[1359:1344] + adder_tree_tier_2_p1_in[1375:1360];
    adder_tree_tier_3_p1_in[703:688] = adder_tree_tier_2_p1_in[1391:1376] + adder_tree_tier_2_p1_in[1407:1392];
    adder_tree_tier_3_p1_in[719:704] = adder_tree_tier_2_p1_in[1423:1408] + adder_tree_tier_2_p1_in[1439:1424];
    adder_tree_tier_3_p1_in[735:720] = adder_tree_tier_2_p1_in[1455:1440] + adder_tree_tier_2_p1_in[1471:1456];
    adder_tree_tier_3_p1_in[751:736] = adder_tree_tier_2_p1_in[1487:1472] + adder_tree_tier_2_p1_in[1503:1488];
    adder_tree_tier_3_p1_in[767:752] = adder_tree_tier_2_p1_in[1519:1504] + adder_tree_tier_2_p1_in[1535:1520];
    adder_tree_tier_3_p1_in[783:768] = adder_tree_tier_2_p1_in[1551:1536] + adder_tree_tier_2_p1_in[1567:1552];
    adder_tree_tier_3_p1_in[799:784] = adder_tree_tier_2_p1_in[1583:1568] + adder_tree_tier_2_p1_in[1599:1584];
    adder_tree_tier_3_p1_in[815:800] = adder_tree_tier_2_p1_in[1615:1600];
    adder_tree_tier_4_p1_in[15:0] = adder_tree_tier_3_p1_in[15:0] + adder_tree_tier_3_p1_in[31:16];
    adder_tree_tier_4_p1_in[31:16] = adder_tree_tier_3_p1_in[47:32] + adder_tree_tier_3_p1_in[63:48];
    adder_tree_tier_4_p1_in[47:32] = adder_tree_tier_3_p1_in[79:64] + adder_tree_tier_3_p1_in[95:80];
    adder_tree_tier_4_p1_in[63:48] = adder_tree_tier_3_p1_in[111:96] + adder_tree_tier_3_p1_in[127:112];
    adder_tree_tier_4_p1_in[79:64] = adder_tree_tier_3_p1_in[143:128] + adder_tree_tier_3_p1_in[159:144];
    adder_tree_tier_4_p1_in[95:80] = adder_tree_tier_3_p1_in[175:160] + adder_tree_tier_3_p1_in[191:176];
    adder_tree_tier_4_p1_in[111:96] = adder_tree_tier_3_p1_in[207:192] + adder_tree_tier_3_p1_in[223:208];
    adder_tree_tier_4_p1_in[127:112] = adder_tree_tier_3_p1_in[239:224] + adder_tree_tier_3_p1_in[255:240];
    adder_tree_tier_4_p1_in[143:128] = adder_tree_tier_3_p1_in[271:256] + adder_tree_tier_3_p1_in[287:272];
    adder_tree_tier_4_p1_in[159:144] = adder_tree_tier_3_p1_in[303:288] + adder_tree_tier_3_p1_in[319:304];
    adder_tree_tier_4_p1_in[175:160] = adder_tree_tier_3_p1_in[335:320] + adder_tree_tier_3_p1_in[351:336];
    adder_tree_tier_4_p1_in[191:176] = adder_tree_tier_3_p1_in[367:352] + adder_tree_tier_3_p1_in[383:368];
    adder_tree_tier_4_p1_in[207:192] = adder_tree_tier_3_p1_in[399:384] + adder_tree_tier_3_p1_in[415:400];
    adder_tree_tier_4_p1_in[223:208] = adder_tree_tier_3_p1_in[431:416] + adder_tree_tier_3_p1_in[447:432];
    adder_tree_tier_4_p1_in[239:224] = adder_tree_tier_3_p1_in[463:448] + adder_tree_tier_3_p1_in[479:464];
    adder_tree_tier_4_p1_in[255:240] = adder_tree_tier_3_p1_in[495:480] + adder_tree_tier_3_p1_in[511:496];
    adder_tree_tier_4_p1_in[271:256] = adder_tree_tier_3_p1_in[527:512] + adder_tree_tier_3_p1_in[543:528];
    adder_tree_tier_4_p1_in[287:272] = adder_tree_tier_3_p1_in[559:544] + adder_tree_tier_3_p1_in[575:560];
    adder_tree_tier_4_p1_in[303:288] = adder_tree_tier_3_p1_in[591:576] + adder_tree_tier_3_p1_in[607:592];
    adder_tree_tier_4_p1_in[319:304] = adder_tree_tier_3_p1_in[623:608] + adder_tree_tier_3_p1_in[639:624];
    adder_tree_tier_4_p1_in[335:320] = adder_tree_tier_3_p1_in[655:640] + adder_tree_tier_3_p1_in[671:656];
    adder_tree_tier_4_p1_in[351:336] = adder_tree_tier_3_p1_in[687:672] + adder_tree_tier_3_p1_in[703:688];
    adder_tree_tier_4_p1_in[367:352] = adder_tree_tier_3_p1_in[719:704] + adder_tree_tier_3_p1_in[735:720];
    adder_tree_tier_4_p1_in[383:368] = adder_tree_tier_3_p1_in[751:736] + adder_tree_tier_3_p1_in[767:752];
    adder_tree_tier_4_p1_in[399:384] = adder_tree_tier_3_p1_in[783:768] + adder_tree_tier_3_p1_in[799:784];
    adder_tree_tier_4_p1_in[415:400] = adder_tree_tier_3_p1_in[815:800];
    adder_tree_tier_5_p1_in[15:0] = adder_tree_tier_4_p1_in[15:0] + adder_tree_tier_4_p1_in[31:16];
    adder_tree_tier_5_p1_in[31:16] = adder_tree_tier_4_p1_in[47:32] + adder_tree_tier_4_p1_in[63:48];
    adder_tree_tier_5_p1_in[47:32] = adder_tree_tier_4_p1_in[79:64] + adder_tree_tier_4_p1_in[95:80];
    adder_tree_tier_5_p1_in[63:48] = adder_tree_tier_4_p1_in[111:96] + adder_tree_tier_4_p1_in[127:112];
    adder_tree_tier_5_p1_in[79:64] = adder_tree_tier_4_p1_in[143:128] + adder_tree_tier_4_p1_in[159:144];
    adder_tree_tier_5_p1_in[95:80] = adder_tree_tier_4_p1_in[175:160] + adder_tree_tier_4_p1_in[191:176];
    adder_tree_tier_5_p1_in[111:96] = adder_tree_tier_4_p1_in[207:192] + adder_tree_tier_4_p1_in[223:208];
    adder_tree_tier_5_p1_in[127:112] = adder_tree_tier_4_p1_in[239:224] + adder_tree_tier_4_p1_in[255:240];
    adder_tree_tier_5_p1_in[143:128] = adder_tree_tier_4_p1_in[271:256] + adder_tree_tier_4_p1_in[287:272];
    adder_tree_tier_5_p1_in[159:144] = adder_tree_tier_4_p1_in[303:288] + adder_tree_tier_4_p1_in[319:304];
    adder_tree_tier_5_p1_in[175:160] = adder_tree_tier_4_p1_in[335:320] + adder_tree_tier_4_p1_in[351:336];
    adder_tree_tier_5_p1_in[191:176] = adder_tree_tier_4_p1_in[367:352] + adder_tree_tier_4_p1_in[383:368];
    adder_tree_tier_5_p1_in[207:192] = adder_tree_tier_4_p1_in[399:384] + adder_tree_tier_4_p1_in[415:400];
    adder_tree_tier_6_p1_in[15:0] = adder_tree_tier_5_p1_in[15:0] + adder_tree_tier_5_p1_in[31:16];
    adder_tree_tier_6_p1_in[31:16] = adder_tree_tier_5_p1_in[47:32] + adder_tree_tier_5_p1_in[63:48];
    adder_tree_tier_6_p1_in[47:32] = adder_tree_tier_5_p1_in[79:64] + adder_tree_tier_5_p1_in[95:80];
    adder_tree_tier_6_p1_in[63:48] = adder_tree_tier_5_p1_in[111:96] + adder_tree_tier_5_p1_in[127:112];
    adder_tree_tier_6_p1_in[79:64] = adder_tree_tier_5_p1_in[143:128] + adder_tree_tier_5_p1_in[159:144];
    adder_tree_tier_6_p1_in[95:80] = adder_tree_tier_5_p1_in[175:160] + adder_tree_tier_5_p1_in[191:176];
    adder_tree_tier_6_p1_in[111:96] = adder_tree_tier_5_p1_in[207:192];
    adder_tree_tier_7_p1_in[15:0] = adder_tree_tier_6_p1_in[15:0] + adder_tree_tier_6_p1_in[31:16];
    adder_tree_tier_7_p1_in[31:16] = adder_tree_tier_6_p1_in[47:32] + adder_tree_tier_6_p1_in[63:48];
    adder_tree_tier_7_p1_in[47:32] = adder_tree_tier_6_p1_in[79:64] + adder_tree_tier_6_p1_in[95:80];
    adder_tree_tier_7_p1_in[63:48] = adder_tree_tier_6_p1_in[111:96];
    adder_tree_tier_8_p1_in[15:0] = adder_tree_tier_7_p1_in[15:0] + adder_tree_tier_7_p1_in[31:16];
    adder_tree_tier_8_p1_in[31:16] = adder_tree_tier_7_p1_in[47:32] + adder_tree_tier_7_p1_in[63:48];
    adder_tree_tier_9_p1_in[15:0] = adder_tree_tier_8_p1_in[15:0] + adder_tree_tier_8_p1_in[31:16];
    val_out_buffer[31:16] = adder_tree_tier_9_p1_in;
  end
  always_ff @(posedge clk or negedge reset) begin
    if (!reset) begin
      history = {(2144){1'b0} };
    end
    else begin
      history = (((history << 32) & {{2112{1'b1}}, {32{1'b0}}}) | cur_val_q);
    end
  end
  assign val_out = val_out_buffer;
endmodule