
module FIR (input logic clk, reset, input logic [15:0] val_in, output logic [15:0] val_out);
  logic [6399:0] history;
  logic [6415:0] value_grid;
  logic [15:0] cur_val_q;
  logic [6415:0] tap_outputs;
  logic [15:0] val_out_buffer;
  assign value_grid = {history, cur_val_q};
  assign cur_val_q = val_in;
  always_comb begin
    logic [6415:0] adder_tree_tier_0_in;
    logic [3215:0] adder_tree_tier_1_in;
    logic [1615:0] adder_tree_tier_2_in;
    logic [815:0] adder_tree_tier_3_in;
    logic [415:0] adder_tree_tier_4_in;
    logic [207:0] adder_tree_tier_5_in;
    logic [111:0] adder_tree_tier_6_in;
    logic [63:0] adder_tree_tier_7_in;
    logic [31:0] adder_tree_tier_8_in;
    logic [15:0] adder_tree_tier_9_in;
    tap_outputs[15:0] = value_grid[15:0] * 11390;
    tap_outputs[31:16] = value_grid[31:16] * 11392;
    tap_outputs[47:32] = value_grid[47:32] * 11391;
    tap_outputs[63:48] = value_grid[63:48] * 11391;
    tap_outputs[79:64] = value_grid[79:64] * 11391;
    tap_outputs[95:80] = value_grid[95:80] * 11390;
    tap_outputs[111:96] = value_grid[111:96] * 11389;
    tap_outputs[127:112] = value_grid[127:112] * 11389;
    tap_outputs[143:128] = value_grid[143:128] * 11389;
    tap_outputs[159:144] = value_grid[159:144] * 11390;
    tap_outputs[175:160] = value_grid[175:160] * 11391;
    tap_outputs[191:176] = value_grid[191:176] * 11392;
    tap_outputs[207:192] = value_grid[207:192] * 11393;
    tap_outputs[223:208] = value_grid[223:208] * 11392;
    tap_outputs[239:224] = value_grid[239:224] * 11390;
    tap_outputs[255:240] = value_grid[255:240] * 11388;
    tap_outputs[271:256] = value_grid[271:256] * 11387;
    tap_outputs[287:272] = value_grid[287:272] * 11387;
    tap_outputs[303:288] = value_grid[303:288] * 11389;
    tap_outputs[319:304] = value_grid[319:304] * 11392;
    tap_outputs[335:320] = value_grid[335:320] * 11394;
    tap_outputs[351:336] = value_grid[351:336] * 11396;
    tap_outputs[367:352] = value_grid[367:352] * 11395;
    tap_outputs[383:368] = value_grid[383:368] * 11391;
    tap_outputs[399:384] = value_grid[399:384] * 11387;
    tap_outputs[415:400] = value_grid[415:400] * 11384;
    tap_outputs[431:416] = value_grid[431:416] * 11383;
    tap_outputs[447:432] = value_grid[447:432] * 11386;
    tap_outputs[463:448] = value_grid[463:448] * 11391;
    tap_outputs[479:464] = value_grid[479:464] * 11397;
    tap_outputs[495:480] = value_grid[495:480] * 11400;
    tap_outputs[511:496] = value_grid[511:496] * 11400;
    tap_outputs[527:512] = value_grid[527:512] * 11395;
    tap_outputs[543:528] = value_grid[543:528] * 11387;
    tap_outputs[559:544] = value_grid[559:544] * 11380;
    tap_outputs[575:560] = value_grid[575:560] * 11377;
    tap_outputs[591:576] = value_grid[591:576] * 11380;
    tap_outputs[607:592] = value_grid[607:592] * 11388;
    tap_outputs[623:608] = value_grid[623:608] * 11399;
    tap_outputs[639:624] = value_grid[639:624] * 11407;
    tap_outputs[655:640] = value_grid[655:640] * 11408;
    tap_outputs[671:656] = value_grid[671:656] * 11401;
    tap_outputs[687:672] = value_grid[687:672] * 11388;
    tap_outputs[703:688] = value_grid[703:688] * 11375;
    tap_outputs[719:704] = value_grid[719:704] * 11367;
    tap_outputs[735:720] = value_grid[735:720] * 11369;
    tap_outputs[751:736] = value_grid[751:736] * 11381;
    tap_outputs[767:752] = value_grid[767:752] * 11399;
    tap_outputs[783:768] = value_grid[783:768] * 11415;
    tap_outputs[799:784] = value_grid[799:784] * 11421;
    tap_outputs[815:800] = value_grid[815:800] * 11413;
    tap_outputs[831:816] = value_grid[831:816] * 11394;
    tap_outputs[847:832] = value_grid[847:832] * 11371;
    tap_outputs[863:848] = value_grid[863:848] * 11355;
    tap_outputs[879:864] = value_grid[879:864] * 11353;
    tap_outputs[895:880] = value_grid[895:880] * 11369;
    tap_outputs[911:896] = value_grid[911:896] * 11396;
    tap_outputs[927:912] = value_grid[927:912] * 11423;
    tap_outputs[943:928] = value_grid[943:928] * 11438;
    tap_outputs[959:944] = value_grid[959:944] * 11433;
    tap_outputs[975:960] = value_grid[975:960] * 11407;
    tap_outputs[991:976] = value_grid[991:976] * 11371;
    tap_outputs[1007:992] = value_grid[1007:992] * 11341;
    tap_outputs[1023:1008] = value_grid[1023:1008] * 11330;
    tap_outputs[1039:1024] = value_grid[1039:1024] * 11347;
    tap_outputs[1055:1040] = value_grid[1055:1040] * 11385;
    tap_outputs[1071:1056] = value_grid[1071:1056] * 11429;
    tap_outputs[1087:1072] = value_grid[1087:1072] * 11460;
    tap_outputs[1103:1088] = value_grid[1103:1088] * 11461;
    tap_outputs[1119:1104] = value_grid[1119:1104] * 11430;
    tap_outputs[1135:1120] = value_grid[1135:1120] * 11378;
    tap_outputs[1151:1136] = value_grid[1151:1136] * 11327;
    tap_outputs[1167:1152] = value_grid[1167:1152] * 11301;
    tap_outputs[1183:1168] = value_grid[1183:1168] * 11314;
    tap_outputs[1199:1184] = value_grid[1199:1184] * 11363;
    tap_outputs[1215:1200] = value_grid[1215:1200] * 11429;
    tap_outputs[1231:1216] = value_grid[1231:1216] * 11483;
    tap_outputs[1247:1232] = value_grid[1247:1232] * 11499;
    tap_outputs[1263:1248] = value_grid[1263:1248] * 11467;
    tap_outputs[1279:1264] = value_grid[1279:1264] * 11396;
    tap_outputs[1295:1280] = value_grid[1295:1280] * 11317;
    tap_outputs[1311:1296] = value_grid[1311:1296] * 11266;
    tap_outputs[1327:1312] = value_grid[1327:1312] * 11267;
    tap_outputs[1343:1328] = value_grid[1343:1328] * 11325;
    tap_outputs[1359:1344] = value_grid[1359:1344] * 11417;
    tap_outputs[1375:1360] = value_grid[1375:1360] * 11505;
    tap_outputs[1391:1376] = value_grid[1391:1376] * 11547;
    tap_outputs[1407:1392] = value_grid[1407:1392] * 11521;
    tap_outputs[1423:1408] = value_grid[1423:1408] * 11433;
    tap_outputs[1439:1424] = value_grid[1439:1424] * 11319;
    tap_outputs[1455:1440] = value_grid[1455:1440] * 11229;
    tap_outputs[1471:1456] = value_grid[1471:1456] * 11206;
    tap_outputs[1487:1472] = value_grid[1487:1472] * 11266;
    tap_outputs[1503:1488] = value_grid[1503:1488] * 11387;
    tap_outputs[1519:1504] = value_grid[1519:1504] * 11519;
    tap_outputs[1535:1520] = value_grid[1535:1520] * 11602;
    tap_outputs[1551:1536] = value_grid[1551:1536] * 11594;
    tap_outputs[1567:1552] = value_grid[1567:1552] * 11493;
    tap_outputs[1583:1568] = value_grid[1583:1568] * 11338;
    tap_outputs[1599:1584] = value_grid[1599:1584] * 11196;
    tap_outputs[1615:1600] = value_grid[1615:1600] * 11132;
    tap_outputs[1631:1616] = value_grid[1631:1616] * 11181;
    tap_outputs[1647:1632] = value_grid[1647:1632] * 11330;
    tap_outputs[1663:1648] = value_grid[1663:1648] * 11516;
    tap_outputs[1679:1664] = value_grid[1679:1664] * 11658;
    tap_outputs[1695:1680] = value_grid[1695:1680] * 11688;
    tap_outputs[1711:1696] = value_grid[1711:1696] * 11584;
    tap_outputs[1727:1712] = value_grid[1727:1712] * 11386;
    tap_outputs[1743:1728] = value_grid[1743:1728] * 11176;
    tap_outputs[1759:1744] = value_grid[1759:1744] * 11049;
    tap_outputs[1775:1760] = value_grid[1775:1760] * 11069;
    tap_outputs[1791:1776] = value_grid[1791:1776] * 11237;
    tap_outputs[1807:1792] = value_grid[1807:1792] * 11485;
    tap_outputs[1823:1808] = value_grid[1823:1808] * 11707;
    tap_outputs[1839:1824] = value_grid[1839:1824] * 11799;
    tap_outputs[1855:1840] = value_grid[1855:1840] * 11712;
    tap_outputs[1871:1856] = value_grid[1871:1856] * 11473;
    tap_outputs[1887:1872] = value_grid[1887:1872] * 11180;
    tap_outputs[1903:1888] = value_grid[1903:1888] * 10965;
    tap_outputs[1919:1904] = value_grid[1919:1904] * 10929;
    tap_outputs[1935:1920] = value_grid[1935:1920] * 11100;
    tap_outputs[1951:1936] = value_grid[1951:1936] * 11414;
    tap_outputs[1967:1952] = value_grid[1967:1952] * 11737;
    tap_outputs[1983:1968] = value_grid[1983:1968] * 11924;
    tap_outputs[1999:1984] = value_grid[1999:1984] * 11880;
    tap_outputs[2015:2000] = value_grid[2015:2000] * 11611;
    tap_outputs[2031:2016] = value_grid[2031:2016] * 11225;
    tap_outputs[2047:2032] = value_grid[2047:2032] * 10891;
    tap_outputs[2063:2048] = value_grid[2063:2048] * 10761;
    tap_outputs[2079:2064] = value_grid[2079:2064] * 10910;
    tap_outputs[2095:2080] = value_grid[2095:2080] * 11285;
    tap_outputs[2111:2096] = value_grid[2111:2096] * 11731;
    tap_outputs[2127:2112] = value_grid[2127:2112] * 12051;
    tap_outputs[2143:2128] = value_grid[2143:2128] * 12090;
    tap_outputs[2159:2144] = value_grid[2159:2144] * 11815;
    tap_outputs[2175:2160] = value_grid[2175:2160] * 11330;
    tap_outputs[2191:2176] = value_grid[2191:2176] * 10842;
    tap_outputs[2207:2192] = value_grid[2207:2192] * 10573;
    tap_outputs[2223:2208] = value_grid[2223:2208] * 10658;
    tap_outputs[2239:2224] = value_grid[2239:2224] * 11080;
    tap_outputs[2255:2240] = value_grid[2255:2240] * 11669;
    tap_outputs[2271:2256] = value_grid[2271:2256] * 12168;
    tap_outputs[2287:2272] = value_grid[2287:2272] * 12345;
    tap_outputs[2303:2288] = value_grid[2303:2288] * 12101;
    tap_outputs[2319:2304] = value_grid[2319:2304] * 11519;
    tap_outputs[2335:2320] = value_grid[2335:2320] * 10842;
    tap_outputs[2351:2336] = value_grid[2351:2336] * 10372;
    tap_outputs[2367:2352] = value_grid[2367:2352] * 10334;
    tap_outputs[2383:2368] = value_grid[2383:2368] * 10773;
    tap_outputs[2399:2384] = value_grid[2399:2384] * 11520;
    tap_outputs[2415:2400] = value_grid[2415:2400] * 12255;
    tap_outputs[2431:2416] = value_grid[2431:2416] * 12645;
    tap_outputs[2447:2432] = value_grid[2447:2432] * 12490;
    tap_outputs[2463:2448] = value_grid[2463:2448] * 11826;
    tap_outputs[2479:2464] = value_grid[2479:2464] * 10921;
    tap_outputs[2495:2480] = value_grid[2495:2480] * 10170;
    tap_outputs[2511:2496] = value_grid[2511:2496] * 9923;
    tap_outputs[2527:2512] = value_grid[2527:2512] * 10327;
    tap_outputs[2543:2528] = value_grid[2543:2528] * 11241;
    tap_outputs[2559:2544] = value_grid[2559:2544] * 12285;
    tap_outputs[2575:2560] = value_grid[2575:2560] * 12995;
    tap_outputs[2591:2576] = value_grid[2591:2576] * 13023;
    tap_outputs[2607:2592] = value_grid[2607:2592] * 12311;
    tap_outputs[2623:2608] = value_grid[2623:2608] * 11128;
    tap_outputs[2639:2624] = value_grid[2639:2624] * 9979;
    tap_outputs[2655:2640] = value_grid[2655:2640] * 9388;
    tap_outputs[2671:2656] = value_grid[2671:2656] * 9667;
    tap_outputs[2687:2672] = value_grid[2687:2672] * 10754;
    tap_outputs[2703:2688] = value_grid[2703:2688] * 12216;
    tap_outputs[2719:2704] = value_grid[2719:2704] * 13416;
    tap_outputs[2735:2720] = value_grid[2735:2720] * 13787;
    tap_outputs[2751:2736] = value_grid[2751:2736] * 13091;
    tap_outputs[2767:2752] = value_grid[2767:2752] * 11557;
    tap_outputs[2783:2768] = value_grid[2783:2768] * 9812;
    tap_outputs[2799:2784] = value_grid[2799:2784] * 8637;
    tap_outputs[2815:2800] = value_grid[2815:2800] * 8619;
    tap_outputs[2831:2816] = value_grid[2831:2816] * 9877;
    tap_outputs[2847:2832] = value_grid[2847:2832] * 11956;
    tap_outputs[2863:2848] = value_grid[2863:2848] * 13985;
    tap_outputs[2879:2864] = value_grid[2879:2864] * 15028;
    tap_outputs[2895:2880] = value_grid[2895:2880] * 14498;
    tap_outputs[2911:2896] = value_grid[2911:2896] * 12463;
    tap_outputs[2927:2912] = value_grid[2927:2912] * 9683;
    tap_outputs[2943:2928] = value_grid[2943:2928] * 7350;
    tap_outputs[2959:2944] = value_grid[2959:2944] * 6602;
    tap_outputs[2975:2960] = value_grid[2975:2960] * 8001;
    tap_outputs[2991:2976] = value_grid[2991:2976] * 11213;
    tap_outputs[3007:2992] = value_grid[3007:2992] * 15026;
    tap_outputs[3023:3008] = value_grid[3023:3008] * 17762;
    tap_outputs[3039:3024] = value_grid[3039:3024] * 17947;
    tap_outputs[3055:3040] = value_grid[3055:3040] * 14992;
    tap_outputs[3071:3056] = value_grid[3071:3056] * 9601;
    tap_outputs[3087:3072] = value_grid[3087:3072] * 3723;
    tap_outputs[3103:3088] = value_grid[3103:3088] * 0;
    tap_outputs[3119:3104] = value_grid[3119:3104] * 874;
    tap_outputs[3135:3120] = value_grid[3135:3120] * 7657;
    tap_outputs[3151:3136] = value_grid[3151:3136] * 19907;
    tap_outputs[3167:3152] = value_grid[3167:3152] * 35362;
    tap_outputs[3183:3168] = value_grid[3183:3168] * 50489;
    tap_outputs[3199:3184] = value_grid[3199:3184] * 61505;
    tap_outputs[3215:3200] = value_grid[3215:3200] * 65535;
    tap_outputs[3231:3216] = value_grid[3231:3216] * 61505;
    tap_outputs[3247:3232] = value_grid[3247:3232] * 50489;
    tap_outputs[3263:3248] = value_grid[3263:3248] * 35362;
    tap_outputs[3279:3264] = value_grid[3279:3264] * 19907;
    tap_outputs[3295:3280] = value_grid[3295:3280] * 7657;
    tap_outputs[3311:3296] = value_grid[3311:3296] * 874;
    tap_outputs[3327:3312] = value_grid[3327:3312] * 0;
    tap_outputs[3343:3328] = value_grid[3343:3328] * 3723;
    tap_outputs[3359:3344] = value_grid[3359:3344] * 9601;
    tap_outputs[3375:3360] = value_grid[3375:3360] * 14992;
    tap_outputs[3391:3376] = value_grid[3391:3376] * 17947;
    tap_outputs[3407:3392] = value_grid[3407:3392] * 17762;
    tap_outputs[3423:3408] = value_grid[3423:3408] * 15026;
    tap_outputs[3439:3424] = value_grid[3439:3424] * 11213;
    tap_outputs[3455:3440] = value_grid[3455:3440] * 8001;
    tap_outputs[3471:3456] = value_grid[3471:3456] * 6602;
    tap_outputs[3487:3472] = value_grid[3487:3472] * 7350;
    tap_outputs[3503:3488] = value_grid[3503:3488] * 9683;
    tap_outputs[3519:3504] = value_grid[3519:3504] * 12463;
    tap_outputs[3535:3520] = value_grid[3535:3520] * 14498;
    tap_outputs[3551:3536] = value_grid[3551:3536] * 15028;
    tap_outputs[3567:3552] = value_grid[3567:3552] * 13985;
    tap_outputs[3583:3568] = value_grid[3583:3568] * 11956;
    tap_outputs[3599:3584] = value_grid[3599:3584] * 9877;
    tap_outputs[3615:3600] = value_grid[3615:3600] * 8619;
    tap_outputs[3631:3616] = value_grid[3631:3616] * 8637;
    tap_outputs[3647:3632] = value_grid[3647:3632] * 9812;
    tap_outputs[3663:3648] = value_grid[3663:3648] * 11557;
    tap_outputs[3679:3664] = value_grid[3679:3664] * 13091;
    tap_outputs[3695:3680] = value_grid[3695:3680] * 13787;
    tap_outputs[3711:3696] = value_grid[3711:3696] * 13416;
    tap_outputs[3727:3712] = value_grid[3727:3712] * 12216;
    tap_outputs[3743:3728] = value_grid[3743:3728] * 10754;
    tap_outputs[3759:3744] = value_grid[3759:3744] * 9667;
    tap_outputs[3775:3760] = value_grid[3775:3760] * 9388;
    tap_outputs[3791:3776] = value_grid[3791:3776] * 9979;
    tap_outputs[3807:3792] = value_grid[3807:3792] * 11128;
    tap_outputs[3823:3808] = value_grid[3823:3808] * 12311;
    tap_outputs[3839:3824] = value_grid[3839:3824] * 13023;
    tap_outputs[3855:3840] = value_grid[3855:3840] * 12995;
    tap_outputs[3871:3856] = value_grid[3871:3856] * 12285;
    tap_outputs[3887:3872] = value_grid[3887:3872] * 11241;
    tap_outputs[3903:3888] = value_grid[3903:3888] * 10327;
    tap_outputs[3919:3904] = value_grid[3919:3904] * 9923;
    tap_outputs[3935:3920] = value_grid[3935:3920] * 10170;
    tap_outputs[3951:3936] = value_grid[3951:3936] * 10921;
    tap_outputs[3967:3952] = value_grid[3967:3952] * 11826;
    tap_outputs[3983:3968] = value_grid[3983:3968] * 12490;
    tap_outputs[3999:3984] = value_grid[3999:3984] * 12645;
    tap_outputs[4015:4000] = value_grid[4015:4000] * 12255;
    tap_outputs[4031:4016] = value_grid[4031:4016] * 11520;
    tap_outputs[4047:4032] = value_grid[4047:4032] * 10773;
    tap_outputs[4063:4048] = value_grid[4063:4048] * 10334;
    tap_outputs[4079:4064] = value_grid[4079:4064] * 10372;
    tap_outputs[4095:4080] = value_grid[4095:4080] * 10842;
    tap_outputs[4111:4096] = value_grid[4111:4096] * 11519;
    tap_outputs[4127:4112] = value_grid[4127:4112] * 12101;
    tap_outputs[4143:4128] = value_grid[4143:4128] * 12345;
    tap_outputs[4159:4144] = value_grid[4159:4144] * 12168;
    tap_outputs[4175:4160] = value_grid[4175:4160] * 11669;
    tap_outputs[4191:4176] = value_grid[4191:4176] * 11080;
    tap_outputs[4207:4192] = value_grid[4207:4192] * 10658;
    tap_outputs[4223:4208] = value_grid[4223:4208] * 10573;
    tap_outputs[4239:4224] = value_grid[4239:4224] * 10842;
    tap_outputs[4255:4240] = value_grid[4255:4240] * 11330;
    tap_outputs[4271:4256] = value_grid[4271:4256] * 11815;
    tap_outputs[4287:4272] = value_grid[4287:4272] * 12090;
    tap_outputs[4303:4288] = value_grid[4303:4288] * 12051;
    tap_outputs[4319:4304] = value_grid[4319:4304] * 11731;
    tap_outputs[4335:4320] = value_grid[4335:4320] * 11285;
    tap_outputs[4351:4336] = value_grid[4351:4336] * 10910;
    tap_outputs[4367:4352] = value_grid[4367:4352] * 10761;
    tap_outputs[4383:4368] = value_grid[4383:4368] * 10891;
    tap_outputs[4399:4384] = value_grid[4399:4384] * 11225;
    tap_outputs[4415:4400] = value_grid[4415:4400] * 11611;
    tap_outputs[4431:4416] = value_grid[4431:4416] * 11880;
    tap_outputs[4447:4432] = value_grid[4447:4432] * 11924;
    tap_outputs[4463:4448] = value_grid[4463:4448] * 11737;
    tap_outputs[4479:4464] = value_grid[4479:4464] * 11414;
    tap_outputs[4495:4480] = value_grid[4495:4480] * 11100;
    tap_outputs[4511:4496] = value_grid[4511:4496] * 10929;
    tap_outputs[4527:4512] = value_grid[4527:4512] * 10965;
    tap_outputs[4543:4528] = value_grid[4543:4528] * 11180;
    tap_outputs[4559:4544] = value_grid[4559:4544] * 11473;
    tap_outputs[4575:4560] = value_grid[4575:4560] * 11712;
    tap_outputs[4591:4576] = value_grid[4591:4576] * 11799;
    tap_outputs[4607:4592] = value_grid[4607:4592] * 11707;
    tap_outputs[4623:4608] = value_grid[4623:4608] * 11485;
    tap_outputs[4639:4624] = value_grid[4639:4624] * 11237;
    tap_outputs[4655:4640] = value_grid[4655:4640] * 11069;
    tap_outputs[4671:4656] = value_grid[4671:4656] * 11049;
    tap_outputs[4687:4672] = value_grid[4687:4672] * 11176;
    tap_outputs[4703:4688] = value_grid[4703:4688] * 11386;
    tap_outputs[4719:4704] = value_grid[4719:4704] * 11584;
    tap_outputs[4735:4720] = value_grid[4735:4720] * 11688;
    tap_outputs[4751:4736] = value_grid[4751:4736] * 11658;
    tap_outputs[4767:4752] = value_grid[4767:4752] * 11516;
    tap_outputs[4783:4768] = value_grid[4783:4768] * 11330;
    tap_outputs[4799:4784] = value_grid[4799:4784] * 11181;
    tap_outputs[4815:4800] = value_grid[4815:4800] * 11132;
    tap_outputs[4831:4816] = value_grid[4831:4816] * 11196;
    tap_outputs[4847:4832] = value_grid[4847:4832] * 11338;
    tap_outputs[4863:4848] = value_grid[4863:4848] * 11493;
    tap_outputs[4879:4864] = value_grid[4879:4864] * 11594;
    tap_outputs[4895:4880] = value_grid[4895:4880] * 11602;
    tap_outputs[4911:4896] = value_grid[4911:4896] * 11519;
    tap_outputs[4927:4912] = value_grid[4927:4912] * 11387;
    tap_outputs[4943:4928] = value_grid[4943:4928] * 11266;
    tap_outputs[4959:4944] = value_grid[4959:4944] * 11206;
    tap_outputs[4975:4960] = value_grid[4975:4960] * 11229;
    tap_outputs[4991:4976] = value_grid[4991:4976] * 11319;
    tap_outputs[5007:4992] = value_grid[5007:4992] * 11433;
    tap_outputs[5023:5008] = value_grid[5023:5008] * 11521;
    tap_outputs[5039:5024] = value_grid[5039:5024] * 11547;
    tap_outputs[5055:5040] = value_grid[5055:5040] * 11505;
    tap_outputs[5071:5056] = value_grid[5071:5056] * 11417;
    tap_outputs[5087:5072] = value_grid[5087:5072] * 11325;
    tap_outputs[5103:5088] = value_grid[5103:5088] * 11267;
    tap_outputs[5119:5104] = value_grid[5119:5104] * 11266;
    tap_outputs[5135:5120] = value_grid[5135:5120] * 11317;
    tap_outputs[5151:5136] = value_grid[5151:5136] * 11396;
    tap_outputs[5167:5152] = value_grid[5167:5152] * 11467;
    tap_outputs[5183:5168] = value_grid[5183:5168] * 11499;
    tap_outputs[5199:5184] = value_grid[5199:5184] * 11483;
    tap_outputs[5215:5200] = value_grid[5215:5200] * 11429;
    tap_outputs[5231:5216] = value_grid[5231:5216] * 11363;
    tap_outputs[5247:5232] = value_grid[5247:5232] * 11314;
    tap_outputs[5263:5248] = value_grid[5263:5248] * 11301;
    tap_outputs[5279:5264] = value_grid[5279:5264] * 11327;
    tap_outputs[5295:5280] = value_grid[5295:5280] * 11378;
    tap_outputs[5311:5296] = value_grid[5311:5296] * 11430;
    tap_outputs[5327:5312] = value_grid[5327:5312] * 11461;
    tap_outputs[5343:5328] = value_grid[5343:5328] * 11460;
    tap_outputs[5359:5344] = value_grid[5359:5344] * 11429;
    tap_outputs[5375:5360] = value_grid[5375:5360] * 11385;
    tap_outputs[5391:5376] = value_grid[5391:5376] * 11347;
    tap_outputs[5407:5392] = value_grid[5407:5392] * 11330;
    tap_outputs[5423:5408] = value_grid[5423:5408] * 11341;
    tap_outputs[5439:5424] = value_grid[5439:5424] * 11371;
    tap_outputs[5455:5440] = value_grid[5455:5440] * 11407;
    tap_outputs[5471:5456] = value_grid[5471:5456] * 11433;
    tap_outputs[5487:5472] = value_grid[5487:5472] * 11438;
    tap_outputs[5503:5488] = value_grid[5503:5488] * 11423;
    tap_outputs[5519:5504] = value_grid[5519:5504] * 11396;
    tap_outputs[5535:5520] = value_grid[5535:5520] * 11369;
    tap_outputs[5551:5536] = value_grid[5551:5536] * 11353;
    tap_outputs[5567:5552] = value_grid[5567:5552] * 11355;
    tap_outputs[5583:5568] = value_grid[5583:5568] * 11371;
    tap_outputs[5599:5584] = value_grid[5599:5584] * 11394;
    tap_outputs[5615:5600] = value_grid[5615:5600] * 11413;
    tap_outputs[5631:5616] = value_grid[5631:5616] * 11421;
    tap_outputs[5647:5632] = value_grid[5647:5632] * 11415;
    tap_outputs[5663:5648] = value_grid[5663:5648] * 11399;
    tap_outputs[5679:5664] = value_grid[5679:5664] * 11381;
    tap_outputs[5695:5680] = value_grid[5695:5680] * 11369;
    tap_outputs[5711:5696] = value_grid[5711:5696] * 11367;
    tap_outputs[5727:5712] = value_grid[5727:5712] * 11375;
    tap_outputs[5743:5728] = value_grid[5743:5728] * 11388;
    tap_outputs[5759:5744] = value_grid[5759:5744] * 11401;
    tap_outputs[5775:5760] = value_grid[5775:5760] * 11408;
    tap_outputs[5791:5776] = value_grid[5791:5776] * 11407;
    tap_outputs[5807:5792] = value_grid[5807:5792] * 11399;
    tap_outputs[5823:5808] = value_grid[5823:5808] * 11388;
    tap_outputs[5839:5824] = value_grid[5839:5824] * 11380;
    tap_outputs[5855:5840] = value_grid[5855:5840] * 11377;
    tap_outputs[5871:5856] = value_grid[5871:5856] * 11380;
    tap_outputs[5887:5872] = value_grid[5887:5872] * 11387;
    tap_outputs[5903:5888] = value_grid[5903:5888] * 11395;
    tap_outputs[5919:5904] = value_grid[5919:5904] * 11400;
    tap_outputs[5935:5920] = value_grid[5935:5920] * 11400;
    tap_outputs[5951:5936] = value_grid[5951:5936] * 11397;
    tap_outputs[5967:5952] = value_grid[5967:5952] * 11391;
    tap_outputs[5983:5968] = value_grid[5983:5968] * 11386;
    tap_outputs[5999:5984] = value_grid[5999:5984] * 11383;
    tap_outputs[6015:6000] = value_grid[6015:6000] * 11384;
    tap_outputs[6031:6016] = value_grid[6031:6016] * 11387;
    tap_outputs[6047:6032] = value_grid[6047:6032] * 11391;
    tap_outputs[6063:6048] = value_grid[6063:6048] * 11395;
    tap_outputs[6079:6064] = value_grid[6079:6064] * 11396;
    tap_outputs[6095:6080] = value_grid[6095:6080] * 11394;
    tap_outputs[6111:6096] = value_grid[6111:6096] * 11392;
    tap_outputs[6127:6112] = value_grid[6127:6112] * 11389;
    tap_outputs[6143:6128] = value_grid[6143:6128] * 11387;
    tap_outputs[6159:6144] = value_grid[6159:6144] * 11387;
    tap_outputs[6175:6160] = value_grid[6175:6160] * 11388;
    tap_outputs[6191:6176] = value_grid[6191:6176] * 11390;
    tap_outputs[6207:6192] = value_grid[6207:6192] * 11392;
    tap_outputs[6223:6208] = value_grid[6223:6208] * 11393;
    tap_outputs[6239:6224] = value_grid[6239:6224] * 11392;
    tap_outputs[6255:6240] = value_grid[6255:6240] * 11391;
    tap_outputs[6271:6256] = value_grid[6271:6256] * 11390;
    tap_outputs[6287:6272] = value_grid[6287:6272] * 11389;
    tap_outputs[6303:6288] = value_grid[6303:6288] * 11389;
    tap_outputs[6319:6304] = value_grid[6319:6304] * 11389;
    tap_outputs[6335:6320] = value_grid[6335:6320] * 11390;
    tap_outputs[6351:6336] = value_grid[6351:6336] * 11391;
    tap_outputs[6367:6352] = value_grid[6367:6352] * 11391;
    tap_outputs[6383:6368] = value_grid[6383:6368] * 11391;
    tap_outputs[6399:6384] = value_grid[6399:6384] * 11392;
    tap_outputs[6415:6400] = value_grid[6415:6400] * 11390;
    adder_tree_tier_0_in = tap_outputs;
    adder_tree_tier_1_in[15:0] = adder_tree_tier_0_in[15:0] + adder_tree_tier_0_in[31:16];
    adder_tree_tier_1_in[31:16] = adder_tree_tier_0_in[47:32] + adder_tree_tier_0_in[63:48];
    adder_tree_tier_1_in[47:32] = adder_tree_tier_0_in[79:64] + adder_tree_tier_0_in[95:80];
    adder_tree_tier_1_in[63:48] = adder_tree_tier_0_in[111:96] + adder_tree_tier_0_in[127:112];
    adder_tree_tier_1_in[79:64] = adder_tree_tier_0_in[143:128] + adder_tree_tier_0_in[159:144];
    adder_tree_tier_1_in[95:80] = adder_tree_tier_0_in[175:160] + adder_tree_tier_0_in[191:176];
    adder_tree_tier_1_in[111:96] = adder_tree_tier_0_in[207:192] + adder_tree_tier_0_in[223:208];
    adder_tree_tier_1_in[127:112] = adder_tree_tier_0_in[239:224] + adder_tree_tier_0_in[255:240];
    adder_tree_tier_1_in[143:128] = adder_tree_tier_0_in[271:256] + adder_tree_tier_0_in[287:272];
    adder_tree_tier_1_in[159:144] = adder_tree_tier_0_in[303:288] + adder_tree_tier_0_in[319:304];
    adder_tree_tier_1_in[175:160] = adder_tree_tier_0_in[335:320] + adder_tree_tier_0_in[351:336];
    adder_tree_tier_1_in[191:176] = adder_tree_tier_0_in[367:352] + adder_tree_tier_0_in[383:368];
    adder_tree_tier_1_in[207:192] = adder_tree_tier_0_in[399:384] + adder_tree_tier_0_in[415:400];
    adder_tree_tier_1_in[223:208] = adder_tree_tier_0_in[431:416] + adder_tree_tier_0_in[447:432];
    adder_tree_tier_1_in[239:224] = adder_tree_tier_0_in[463:448] + adder_tree_tier_0_in[479:464];
    adder_tree_tier_1_in[255:240] = adder_tree_tier_0_in[495:480] + adder_tree_tier_0_in[511:496];
    adder_tree_tier_1_in[271:256] = adder_tree_tier_0_in[527:512] + adder_tree_tier_0_in[543:528];
    adder_tree_tier_1_in[287:272] = adder_tree_tier_0_in[559:544] + adder_tree_tier_0_in[575:560];
    adder_tree_tier_1_in[303:288] = adder_tree_tier_0_in[591:576] + adder_tree_tier_0_in[607:592];
    adder_tree_tier_1_in[319:304] = adder_tree_tier_0_in[623:608] + adder_tree_tier_0_in[639:624];
    adder_tree_tier_1_in[335:320] = adder_tree_tier_0_in[655:640] + adder_tree_tier_0_in[671:656];
    adder_tree_tier_1_in[351:336] = adder_tree_tier_0_in[687:672] + adder_tree_tier_0_in[703:688];
    adder_tree_tier_1_in[367:352] = adder_tree_tier_0_in[719:704] + adder_tree_tier_0_in[735:720];
    adder_tree_tier_1_in[383:368] = adder_tree_tier_0_in[751:736] + adder_tree_tier_0_in[767:752];
    adder_tree_tier_1_in[399:384] = adder_tree_tier_0_in[783:768] + adder_tree_tier_0_in[799:784];
    adder_tree_tier_1_in[415:400] = adder_tree_tier_0_in[815:800] + adder_tree_tier_0_in[831:816];
    adder_tree_tier_1_in[431:416] = adder_tree_tier_0_in[847:832] + adder_tree_tier_0_in[863:848];
    adder_tree_tier_1_in[447:432] = adder_tree_tier_0_in[879:864] + adder_tree_tier_0_in[895:880];
    adder_tree_tier_1_in[463:448] = adder_tree_tier_0_in[911:896] + adder_tree_tier_0_in[927:912];
    adder_tree_tier_1_in[479:464] = adder_tree_tier_0_in[943:928] + adder_tree_tier_0_in[959:944];
    adder_tree_tier_1_in[495:480] = adder_tree_tier_0_in[975:960] + adder_tree_tier_0_in[991:976];
    adder_tree_tier_1_in[511:496] = adder_tree_tier_0_in[1007:992] + adder_tree_tier_0_in[1023:1008];
    adder_tree_tier_1_in[527:512] = adder_tree_tier_0_in[1039:1024] + adder_tree_tier_0_in[1055:1040];
    adder_tree_tier_1_in[543:528] = adder_tree_tier_0_in[1071:1056] + adder_tree_tier_0_in[1087:1072];
    adder_tree_tier_1_in[559:544] = adder_tree_tier_0_in[1103:1088] + adder_tree_tier_0_in[1119:1104];
    adder_tree_tier_1_in[575:560] = adder_tree_tier_0_in[1135:1120] + adder_tree_tier_0_in[1151:1136];
    adder_tree_tier_1_in[591:576] = adder_tree_tier_0_in[1167:1152] + adder_tree_tier_0_in[1183:1168];
    adder_tree_tier_1_in[607:592] = adder_tree_tier_0_in[1199:1184] + adder_tree_tier_0_in[1215:1200];
    adder_tree_tier_1_in[623:608] = adder_tree_tier_0_in[1231:1216] + adder_tree_tier_0_in[1247:1232];
    adder_tree_tier_1_in[639:624] = adder_tree_tier_0_in[1263:1248] + adder_tree_tier_0_in[1279:1264];
    adder_tree_tier_1_in[655:640] = adder_tree_tier_0_in[1295:1280] + adder_tree_tier_0_in[1311:1296];
    adder_tree_tier_1_in[671:656] = adder_tree_tier_0_in[1327:1312] + adder_tree_tier_0_in[1343:1328];
    adder_tree_tier_1_in[687:672] = adder_tree_tier_0_in[1359:1344] + adder_tree_tier_0_in[1375:1360];
    adder_tree_tier_1_in[703:688] = adder_tree_tier_0_in[1391:1376] + adder_tree_tier_0_in[1407:1392];
    adder_tree_tier_1_in[719:704] = adder_tree_tier_0_in[1423:1408] + adder_tree_tier_0_in[1439:1424];
    adder_tree_tier_1_in[735:720] = adder_tree_tier_0_in[1455:1440] + adder_tree_tier_0_in[1471:1456];
    adder_tree_tier_1_in[751:736] = adder_tree_tier_0_in[1487:1472] + adder_tree_tier_0_in[1503:1488];
    adder_tree_tier_1_in[767:752] = adder_tree_tier_0_in[1519:1504] + adder_tree_tier_0_in[1535:1520];
    adder_tree_tier_1_in[783:768] = adder_tree_tier_0_in[1551:1536] + adder_tree_tier_0_in[1567:1552];
    adder_tree_tier_1_in[799:784] = adder_tree_tier_0_in[1583:1568] + adder_tree_tier_0_in[1599:1584];
    adder_tree_tier_1_in[815:800] = adder_tree_tier_0_in[1615:1600] + adder_tree_tier_0_in[1631:1616];
    adder_tree_tier_1_in[831:816] = adder_tree_tier_0_in[1647:1632] + adder_tree_tier_0_in[1663:1648];
    adder_tree_tier_1_in[847:832] = adder_tree_tier_0_in[1679:1664] + adder_tree_tier_0_in[1695:1680];
    adder_tree_tier_1_in[863:848] = adder_tree_tier_0_in[1711:1696] + adder_tree_tier_0_in[1727:1712];
    adder_tree_tier_1_in[879:864] = adder_tree_tier_0_in[1743:1728] + adder_tree_tier_0_in[1759:1744];
    adder_tree_tier_1_in[895:880] = adder_tree_tier_0_in[1775:1760] + adder_tree_tier_0_in[1791:1776];
    adder_tree_tier_1_in[911:896] = adder_tree_tier_0_in[1807:1792] + adder_tree_tier_0_in[1823:1808];
    adder_tree_tier_1_in[927:912] = adder_tree_tier_0_in[1839:1824] + adder_tree_tier_0_in[1855:1840];
    adder_tree_tier_1_in[943:928] = adder_tree_tier_0_in[1871:1856] + adder_tree_tier_0_in[1887:1872];
    adder_tree_tier_1_in[959:944] = adder_tree_tier_0_in[1903:1888] + adder_tree_tier_0_in[1919:1904];
    adder_tree_tier_1_in[975:960] = adder_tree_tier_0_in[1935:1920] + adder_tree_tier_0_in[1951:1936];
    adder_tree_tier_1_in[991:976] = adder_tree_tier_0_in[1967:1952] + adder_tree_tier_0_in[1983:1968];
    adder_tree_tier_1_in[1007:992] = adder_tree_tier_0_in[1999:1984] + adder_tree_tier_0_in[2015:2000];
    adder_tree_tier_1_in[1023:1008] = adder_tree_tier_0_in[2031:2016] + adder_tree_tier_0_in[2047:2032];
    adder_tree_tier_1_in[1039:1024] = adder_tree_tier_0_in[2063:2048] + adder_tree_tier_0_in[2079:2064];
    adder_tree_tier_1_in[1055:1040] = adder_tree_tier_0_in[2095:2080] + adder_tree_tier_0_in[2111:2096];
    adder_tree_tier_1_in[1071:1056] = adder_tree_tier_0_in[2127:2112] + adder_tree_tier_0_in[2143:2128];
    adder_tree_tier_1_in[1087:1072] = adder_tree_tier_0_in[2159:2144] + adder_tree_tier_0_in[2175:2160];
    adder_tree_tier_1_in[1103:1088] = adder_tree_tier_0_in[2191:2176] + adder_tree_tier_0_in[2207:2192];
    adder_tree_tier_1_in[1119:1104] = adder_tree_tier_0_in[2223:2208] + adder_tree_tier_0_in[2239:2224];
    adder_tree_tier_1_in[1135:1120] = adder_tree_tier_0_in[2255:2240] + adder_tree_tier_0_in[2271:2256];
    adder_tree_tier_1_in[1151:1136] = adder_tree_tier_0_in[2287:2272] + adder_tree_tier_0_in[2303:2288];
    adder_tree_tier_1_in[1167:1152] = adder_tree_tier_0_in[2319:2304] + adder_tree_tier_0_in[2335:2320];
    adder_tree_tier_1_in[1183:1168] = adder_tree_tier_0_in[2351:2336] + adder_tree_tier_0_in[2367:2352];
    adder_tree_tier_1_in[1199:1184] = adder_tree_tier_0_in[2383:2368] + adder_tree_tier_0_in[2399:2384];
    adder_tree_tier_1_in[1215:1200] = adder_tree_tier_0_in[2415:2400] + adder_tree_tier_0_in[2431:2416];
    adder_tree_tier_1_in[1231:1216] = adder_tree_tier_0_in[2447:2432] + adder_tree_tier_0_in[2463:2448];
    adder_tree_tier_1_in[1247:1232] = adder_tree_tier_0_in[2479:2464] + adder_tree_tier_0_in[2495:2480];
    adder_tree_tier_1_in[1263:1248] = adder_tree_tier_0_in[2511:2496] + adder_tree_tier_0_in[2527:2512];
    adder_tree_tier_1_in[1279:1264] = adder_tree_tier_0_in[2543:2528] + adder_tree_tier_0_in[2559:2544];
    adder_tree_tier_1_in[1295:1280] = adder_tree_tier_0_in[2575:2560] + adder_tree_tier_0_in[2591:2576];
    adder_tree_tier_1_in[1311:1296] = adder_tree_tier_0_in[2607:2592] + adder_tree_tier_0_in[2623:2608];
    adder_tree_tier_1_in[1327:1312] = adder_tree_tier_0_in[2639:2624] + adder_tree_tier_0_in[2655:2640];
    adder_tree_tier_1_in[1343:1328] = adder_tree_tier_0_in[2671:2656] + adder_tree_tier_0_in[2687:2672];
    adder_tree_tier_1_in[1359:1344] = adder_tree_tier_0_in[2703:2688] + adder_tree_tier_0_in[2719:2704];
    adder_tree_tier_1_in[1375:1360] = adder_tree_tier_0_in[2735:2720] + adder_tree_tier_0_in[2751:2736];
    adder_tree_tier_1_in[1391:1376] = adder_tree_tier_0_in[2767:2752] + adder_tree_tier_0_in[2783:2768];
    adder_tree_tier_1_in[1407:1392] = adder_tree_tier_0_in[2799:2784] + adder_tree_tier_0_in[2815:2800];
    adder_tree_tier_1_in[1423:1408] = adder_tree_tier_0_in[2831:2816] + adder_tree_tier_0_in[2847:2832];
    adder_tree_tier_1_in[1439:1424] = adder_tree_tier_0_in[2863:2848] + adder_tree_tier_0_in[2879:2864];
    adder_tree_tier_1_in[1455:1440] = adder_tree_tier_0_in[2895:2880] + adder_tree_tier_0_in[2911:2896];
    adder_tree_tier_1_in[1471:1456] = adder_tree_tier_0_in[2927:2912] + adder_tree_tier_0_in[2943:2928];
    adder_tree_tier_1_in[1487:1472] = adder_tree_tier_0_in[2959:2944] + adder_tree_tier_0_in[2975:2960];
    adder_tree_tier_1_in[1503:1488] = adder_tree_tier_0_in[2991:2976] + adder_tree_tier_0_in[3007:2992];
    adder_tree_tier_1_in[1519:1504] = adder_tree_tier_0_in[3023:3008] + adder_tree_tier_0_in[3039:3024];
    adder_tree_tier_1_in[1535:1520] = adder_tree_tier_0_in[3055:3040] + adder_tree_tier_0_in[3071:3056];
    adder_tree_tier_1_in[1551:1536] = adder_tree_tier_0_in[3087:3072] + adder_tree_tier_0_in[3103:3088];
    adder_tree_tier_1_in[1567:1552] = adder_tree_tier_0_in[3119:3104] + adder_tree_tier_0_in[3135:3120];
    adder_tree_tier_1_in[1583:1568] = adder_tree_tier_0_in[3151:3136] + adder_tree_tier_0_in[3167:3152];
    adder_tree_tier_1_in[1599:1584] = adder_tree_tier_0_in[3183:3168] + adder_tree_tier_0_in[3199:3184];
    adder_tree_tier_1_in[1615:1600] = adder_tree_tier_0_in[3215:3200] + adder_tree_tier_0_in[3231:3216];
    adder_tree_tier_1_in[1631:1616] = adder_tree_tier_0_in[3247:3232] + adder_tree_tier_0_in[3263:3248];
    adder_tree_tier_1_in[1647:1632] = adder_tree_tier_0_in[3279:3264] + adder_tree_tier_0_in[3295:3280];
    adder_tree_tier_1_in[1663:1648] = adder_tree_tier_0_in[3311:3296] + adder_tree_tier_0_in[3327:3312];
    adder_tree_tier_1_in[1679:1664] = adder_tree_tier_0_in[3343:3328] + adder_tree_tier_0_in[3359:3344];
    adder_tree_tier_1_in[1695:1680] = adder_tree_tier_0_in[3375:3360] + adder_tree_tier_0_in[3391:3376];
    adder_tree_tier_1_in[1711:1696] = adder_tree_tier_0_in[3407:3392] + adder_tree_tier_0_in[3423:3408];
    adder_tree_tier_1_in[1727:1712] = adder_tree_tier_0_in[3439:3424] + adder_tree_tier_0_in[3455:3440];
    adder_tree_tier_1_in[1743:1728] = adder_tree_tier_0_in[3471:3456] + adder_tree_tier_0_in[3487:3472];
    adder_tree_tier_1_in[1759:1744] = adder_tree_tier_0_in[3503:3488] + adder_tree_tier_0_in[3519:3504];
    adder_tree_tier_1_in[1775:1760] = adder_tree_tier_0_in[3535:3520] + adder_tree_tier_0_in[3551:3536];
    adder_tree_tier_1_in[1791:1776] = adder_tree_tier_0_in[3567:3552] + adder_tree_tier_0_in[3583:3568];
    adder_tree_tier_1_in[1807:1792] = adder_tree_tier_0_in[3599:3584] + adder_tree_tier_0_in[3615:3600];
    adder_tree_tier_1_in[1823:1808] = adder_tree_tier_0_in[3631:3616] + adder_tree_tier_0_in[3647:3632];
    adder_tree_tier_1_in[1839:1824] = adder_tree_tier_0_in[3663:3648] + adder_tree_tier_0_in[3679:3664];
    adder_tree_tier_1_in[1855:1840] = adder_tree_tier_0_in[3695:3680] + adder_tree_tier_0_in[3711:3696];
    adder_tree_tier_1_in[1871:1856] = adder_tree_tier_0_in[3727:3712] + adder_tree_tier_0_in[3743:3728];
    adder_tree_tier_1_in[1887:1872] = adder_tree_tier_0_in[3759:3744] + adder_tree_tier_0_in[3775:3760];
    adder_tree_tier_1_in[1903:1888] = adder_tree_tier_0_in[3791:3776] + adder_tree_tier_0_in[3807:3792];
    adder_tree_tier_1_in[1919:1904] = adder_tree_tier_0_in[3823:3808] + adder_tree_tier_0_in[3839:3824];
    adder_tree_tier_1_in[1935:1920] = adder_tree_tier_0_in[3855:3840] + adder_tree_tier_0_in[3871:3856];
    adder_tree_tier_1_in[1951:1936] = adder_tree_tier_0_in[3887:3872] + adder_tree_tier_0_in[3903:3888];
    adder_tree_tier_1_in[1967:1952] = adder_tree_tier_0_in[3919:3904] + adder_tree_tier_0_in[3935:3920];
    adder_tree_tier_1_in[1983:1968] = adder_tree_tier_0_in[3951:3936] + adder_tree_tier_0_in[3967:3952];
    adder_tree_tier_1_in[1999:1984] = adder_tree_tier_0_in[3983:3968] + adder_tree_tier_0_in[3999:3984];
    adder_tree_tier_1_in[2015:2000] = adder_tree_tier_0_in[4015:4000] + adder_tree_tier_0_in[4031:4016];
    adder_tree_tier_1_in[2031:2016] = adder_tree_tier_0_in[4047:4032] + adder_tree_tier_0_in[4063:4048];
    adder_tree_tier_1_in[2047:2032] = adder_tree_tier_0_in[4079:4064] + adder_tree_tier_0_in[4095:4080];
    adder_tree_tier_1_in[2063:2048] = adder_tree_tier_0_in[4111:4096] + adder_tree_tier_0_in[4127:4112];
    adder_tree_tier_1_in[2079:2064] = adder_tree_tier_0_in[4143:4128] + adder_tree_tier_0_in[4159:4144];
    adder_tree_tier_1_in[2095:2080] = adder_tree_tier_0_in[4175:4160] + adder_tree_tier_0_in[4191:4176];
    adder_tree_tier_1_in[2111:2096] = adder_tree_tier_0_in[4207:4192] + adder_tree_tier_0_in[4223:4208];
    adder_tree_tier_1_in[2127:2112] = adder_tree_tier_0_in[4239:4224] + adder_tree_tier_0_in[4255:4240];
    adder_tree_tier_1_in[2143:2128] = adder_tree_tier_0_in[4271:4256] + adder_tree_tier_0_in[4287:4272];
    adder_tree_tier_1_in[2159:2144] = adder_tree_tier_0_in[4303:4288] + adder_tree_tier_0_in[4319:4304];
    adder_tree_tier_1_in[2175:2160] = adder_tree_tier_0_in[4335:4320] + adder_tree_tier_0_in[4351:4336];
    adder_tree_tier_1_in[2191:2176] = adder_tree_tier_0_in[4367:4352] + adder_tree_tier_0_in[4383:4368];
    adder_tree_tier_1_in[2207:2192] = adder_tree_tier_0_in[4399:4384] + adder_tree_tier_0_in[4415:4400];
    adder_tree_tier_1_in[2223:2208] = adder_tree_tier_0_in[4431:4416] + adder_tree_tier_0_in[4447:4432];
    adder_tree_tier_1_in[2239:2224] = adder_tree_tier_0_in[4463:4448] + adder_tree_tier_0_in[4479:4464];
    adder_tree_tier_1_in[2255:2240] = adder_tree_tier_0_in[4495:4480] + adder_tree_tier_0_in[4511:4496];
    adder_tree_tier_1_in[2271:2256] = adder_tree_tier_0_in[4527:4512] + adder_tree_tier_0_in[4543:4528];
    adder_tree_tier_1_in[2287:2272] = adder_tree_tier_0_in[4559:4544] + adder_tree_tier_0_in[4575:4560];
    adder_tree_tier_1_in[2303:2288] = adder_tree_tier_0_in[4591:4576] + adder_tree_tier_0_in[4607:4592];
    adder_tree_tier_1_in[2319:2304] = adder_tree_tier_0_in[4623:4608] + adder_tree_tier_0_in[4639:4624];
    adder_tree_tier_1_in[2335:2320] = adder_tree_tier_0_in[4655:4640] + adder_tree_tier_0_in[4671:4656];
    adder_tree_tier_1_in[2351:2336] = adder_tree_tier_0_in[4687:4672] + adder_tree_tier_0_in[4703:4688];
    adder_tree_tier_1_in[2367:2352] = adder_tree_tier_0_in[4719:4704] + adder_tree_tier_0_in[4735:4720];
    adder_tree_tier_1_in[2383:2368] = adder_tree_tier_0_in[4751:4736] + adder_tree_tier_0_in[4767:4752];
    adder_tree_tier_1_in[2399:2384] = adder_tree_tier_0_in[4783:4768] + adder_tree_tier_0_in[4799:4784];
    adder_tree_tier_1_in[2415:2400] = adder_tree_tier_0_in[4815:4800] + adder_tree_tier_0_in[4831:4816];
    adder_tree_tier_1_in[2431:2416] = adder_tree_tier_0_in[4847:4832] + adder_tree_tier_0_in[4863:4848];
    adder_tree_tier_1_in[2447:2432] = adder_tree_tier_0_in[4879:4864] + adder_tree_tier_0_in[4895:4880];
    adder_tree_tier_1_in[2463:2448] = adder_tree_tier_0_in[4911:4896] + adder_tree_tier_0_in[4927:4912];
    adder_tree_tier_1_in[2479:2464] = adder_tree_tier_0_in[4943:4928] + adder_tree_tier_0_in[4959:4944];
    adder_tree_tier_1_in[2495:2480] = adder_tree_tier_0_in[4975:4960] + adder_tree_tier_0_in[4991:4976];
    adder_tree_tier_1_in[2511:2496] = adder_tree_tier_0_in[5007:4992] + adder_tree_tier_0_in[5023:5008];
    adder_tree_tier_1_in[2527:2512] = adder_tree_tier_0_in[5039:5024] + adder_tree_tier_0_in[5055:5040];
    adder_tree_tier_1_in[2543:2528] = adder_tree_tier_0_in[5071:5056] + adder_tree_tier_0_in[5087:5072];
    adder_tree_tier_1_in[2559:2544] = adder_tree_tier_0_in[5103:5088] + adder_tree_tier_0_in[5119:5104];
    adder_tree_tier_1_in[2575:2560] = adder_tree_tier_0_in[5135:5120] + adder_tree_tier_0_in[5151:5136];
    adder_tree_tier_1_in[2591:2576] = adder_tree_tier_0_in[5167:5152] + adder_tree_tier_0_in[5183:5168];
    adder_tree_tier_1_in[2607:2592] = adder_tree_tier_0_in[5199:5184] + adder_tree_tier_0_in[5215:5200];
    adder_tree_tier_1_in[2623:2608] = adder_tree_tier_0_in[5231:5216] + adder_tree_tier_0_in[5247:5232];
    adder_tree_tier_1_in[2639:2624] = adder_tree_tier_0_in[5263:5248] + adder_tree_tier_0_in[5279:5264];
    adder_tree_tier_1_in[2655:2640] = adder_tree_tier_0_in[5295:5280] + adder_tree_tier_0_in[5311:5296];
    adder_tree_tier_1_in[2671:2656] = adder_tree_tier_0_in[5327:5312] + adder_tree_tier_0_in[5343:5328];
    adder_tree_tier_1_in[2687:2672] = adder_tree_tier_0_in[5359:5344] + adder_tree_tier_0_in[5375:5360];
    adder_tree_tier_1_in[2703:2688] = adder_tree_tier_0_in[5391:5376] + adder_tree_tier_0_in[5407:5392];
    adder_tree_tier_1_in[2719:2704] = adder_tree_tier_0_in[5423:5408] + adder_tree_tier_0_in[5439:5424];
    adder_tree_tier_1_in[2735:2720] = adder_tree_tier_0_in[5455:5440] + adder_tree_tier_0_in[5471:5456];
    adder_tree_tier_1_in[2751:2736] = adder_tree_tier_0_in[5487:5472] + adder_tree_tier_0_in[5503:5488];
    adder_tree_tier_1_in[2767:2752] = adder_tree_tier_0_in[5519:5504] + adder_tree_tier_0_in[5535:5520];
    adder_tree_tier_1_in[2783:2768] = adder_tree_tier_0_in[5551:5536] + adder_tree_tier_0_in[5567:5552];
    adder_tree_tier_1_in[2799:2784] = adder_tree_tier_0_in[5583:5568] + adder_tree_tier_0_in[5599:5584];
    adder_tree_tier_1_in[2815:2800] = adder_tree_tier_0_in[5615:5600] + adder_tree_tier_0_in[5631:5616];
    adder_tree_tier_1_in[2831:2816] = adder_tree_tier_0_in[5647:5632] + adder_tree_tier_0_in[5663:5648];
    adder_tree_tier_1_in[2847:2832] = adder_tree_tier_0_in[5679:5664] + adder_tree_tier_0_in[5695:5680];
    adder_tree_tier_1_in[2863:2848] = adder_tree_tier_0_in[5711:5696] + adder_tree_tier_0_in[5727:5712];
    adder_tree_tier_1_in[2879:2864] = adder_tree_tier_0_in[5743:5728] + adder_tree_tier_0_in[5759:5744];
    adder_tree_tier_1_in[2895:2880] = adder_tree_tier_0_in[5775:5760] + adder_tree_tier_0_in[5791:5776];
    adder_tree_tier_1_in[2911:2896] = adder_tree_tier_0_in[5807:5792] + adder_tree_tier_0_in[5823:5808];
    adder_tree_tier_1_in[2927:2912] = adder_tree_tier_0_in[5839:5824] + adder_tree_tier_0_in[5855:5840];
    adder_tree_tier_1_in[2943:2928] = adder_tree_tier_0_in[5871:5856] + adder_tree_tier_0_in[5887:5872];
    adder_tree_tier_1_in[2959:2944] = adder_tree_tier_0_in[5903:5888] + adder_tree_tier_0_in[5919:5904];
    adder_tree_tier_1_in[2975:2960] = adder_tree_tier_0_in[5935:5920] + adder_tree_tier_0_in[5951:5936];
    adder_tree_tier_1_in[2991:2976] = adder_tree_tier_0_in[5967:5952] + adder_tree_tier_0_in[5983:5968];
    adder_tree_tier_1_in[3007:2992] = adder_tree_tier_0_in[5999:5984] + adder_tree_tier_0_in[6015:6000];
    adder_tree_tier_1_in[3023:3008] = adder_tree_tier_0_in[6031:6016] + adder_tree_tier_0_in[6047:6032];
    adder_tree_tier_1_in[3039:3024] = adder_tree_tier_0_in[6063:6048] + adder_tree_tier_0_in[6079:6064];
    adder_tree_tier_1_in[3055:3040] = adder_tree_tier_0_in[6095:6080] + adder_tree_tier_0_in[6111:6096];
    adder_tree_tier_1_in[3071:3056] = adder_tree_tier_0_in[6127:6112] + adder_tree_tier_0_in[6143:6128];
    adder_tree_tier_1_in[3087:3072] = adder_tree_tier_0_in[6159:6144] + adder_tree_tier_0_in[6175:6160];
    adder_tree_tier_1_in[3103:3088] = adder_tree_tier_0_in[6191:6176] + adder_tree_tier_0_in[6207:6192];
    adder_tree_tier_1_in[3119:3104] = adder_tree_tier_0_in[6223:6208] + adder_tree_tier_0_in[6239:6224];
    adder_tree_tier_1_in[3135:3120] = adder_tree_tier_0_in[6255:6240] + adder_tree_tier_0_in[6271:6256];
    adder_tree_tier_1_in[3151:3136] = adder_tree_tier_0_in[6287:6272] + adder_tree_tier_0_in[6303:6288];
    adder_tree_tier_1_in[3167:3152] = adder_tree_tier_0_in[6319:6304] + adder_tree_tier_0_in[6335:6320];
    adder_tree_tier_1_in[3183:3168] = adder_tree_tier_0_in[6351:6336] + adder_tree_tier_0_in[6367:6352];
    adder_tree_tier_1_in[3199:3184] = adder_tree_tier_0_in[6383:6368] + adder_tree_tier_0_in[6399:6384];
    adder_tree_tier_1_in[3215:3200] = adder_tree_tier_0_in[6415:6400];
    adder_tree_tier_2_in[15:0] = adder_tree_tier_1_in[15:0] + adder_tree_tier_1_in[31:16];
    adder_tree_tier_2_in[31:16] = adder_tree_tier_1_in[47:32] + adder_tree_tier_1_in[63:48];
    adder_tree_tier_2_in[47:32] = adder_tree_tier_1_in[79:64] + adder_tree_tier_1_in[95:80];
    adder_tree_tier_2_in[63:48] = adder_tree_tier_1_in[111:96] + adder_tree_tier_1_in[127:112];
    adder_tree_tier_2_in[79:64] = adder_tree_tier_1_in[143:128] + adder_tree_tier_1_in[159:144];
    adder_tree_tier_2_in[95:80] = adder_tree_tier_1_in[175:160] + adder_tree_tier_1_in[191:176];
    adder_tree_tier_2_in[111:96] = adder_tree_tier_1_in[207:192] + adder_tree_tier_1_in[223:208];
    adder_tree_tier_2_in[127:112] = adder_tree_tier_1_in[239:224] + adder_tree_tier_1_in[255:240];
    adder_tree_tier_2_in[143:128] = adder_tree_tier_1_in[271:256] + adder_tree_tier_1_in[287:272];
    adder_tree_tier_2_in[159:144] = adder_tree_tier_1_in[303:288] + adder_tree_tier_1_in[319:304];
    adder_tree_tier_2_in[175:160] = adder_tree_tier_1_in[335:320] + adder_tree_tier_1_in[351:336];
    adder_tree_tier_2_in[191:176] = adder_tree_tier_1_in[367:352] + adder_tree_tier_1_in[383:368];
    adder_tree_tier_2_in[207:192] = adder_tree_tier_1_in[399:384] + adder_tree_tier_1_in[415:400];
    adder_tree_tier_2_in[223:208] = adder_tree_tier_1_in[431:416] + adder_tree_tier_1_in[447:432];
    adder_tree_tier_2_in[239:224] = adder_tree_tier_1_in[463:448] + adder_tree_tier_1_in[479:464];
    adder_tree_tier_2_in[255:240] = adder_tree_tier_1_in[495:480] + adder_tree_tier_1_in[511:496];
    adder_tree_tier_2_in[271:256] = adder_tree_tier_1_in[527:512] + adder_tree_tier_1_in[543:528];
    adder_tree_tier_2_in[287:272] = adder_tree_tier_1_in[559:544] + adder_tree_tier_1_in[575:560];
    adder_tree_tier_2_in[303:288] = adder_tree_tier_1_in[591:576] + adder_tree_tier_1_in[607:592];
    adder_tree_tier_2_in[319:304] = adder_tree_tier_1_in[623:608] + adder_tree_tier_1_in[639:624];
    adder_tree_tier_2_in[335:320] = adder_tree_tier_1_in[655:640] + adder_tree_tier_1_in[671:656];
    adder_tree_tier_2_in[351:336] = adder_tree_tier_1_in[687:672] + adder_tree_tier_1_in[703:688];
    adder_tree_tier_2_in[367:352] = adder_tree_tier_1_in[719:704] + adder_tree_tier_1_in[735:720];
    adder_tree_tier_2_in[383:368] = adder_tree_tier_1_in[751:736] + adder_tree_tier_1_in[767:752];
    adder_tree_tier_2_in[399:384] = adder_tree_tier_1_in[783:768] + adder_tree_tier_1_in[799:784];
    adder_tree_tier_2_in[415:400] = adder_tree_tier_1_in[815:800] + adder_tree_tier_1_in[831:816];
    adder_tree_tier_2_in[431:416] = adder_tree_tier_1_in[847:832] + adder_tree_tier_1_in[863:848];
    adder_tree_tier_2_in[447:432] = adder_tree_tier_1_in[879:864] + adder_tree_tier_1_in[895:880];
    adder_tree_tier_2_in[463:448] = adder_tree_tier_1_in[911:896] + adder_tree_tier_1_in[927:912];
    adder_tree_tier_2_in[479:464] = adder_tree_tier_1_in[943:928] + adder_tree_tier_1_in[959:944];
    adder_tree_tier_2_in[495:480] = adder_tree_tier_1_in[975:960] + adder_tree_tier_1_in[991:976];
    adder_tree_tier_2_in[511:496] = adder_tree_tier_1_in[1007:992] + adder_tree_tier_1_in[1023:1008];
    adder_tree_tier_2_in[527:512] = adder_tree_tier_1_in[1039:1024] + adder_tree_tier_1_in[1055:1040];
    adder_tree_tier_2_in[543:528] = adder_tree_tier_1_in[1071:1056] + adder_tree_tier_1_in[1087:1072];
    adder_tree_tier_2_in[559:544] = adder_tree_tier_1_in[1103:1088] + adder_tree_tier_1_in[1119:1104];
    adder_tree_tier_2_in[575:560] = adder_tree_tier_1_in[1135:1120] + adder_tree_tier_1_in[1151:1136];
    adder_tree_tier_2_in[591:576] = adder_tree_tier_1_in[1167:1152] + adder_tree_tier_1_in[1183:1168];
    adder_tree_tier_2_in[607:592] = adder_tree_tier_1_in[1199:1184] + adder_tree_tier_1_in[1215:1200];
    adder_tree_tier_2_in[623:608] = adder_tree_tier_1_in[1231:1216] + adder_tree_tier_1_in[1247:1232];
    adder_tree_tier_2_in[639:624] = adder_tree_tier_1_in[1263:1248] + adder_tree_tier_1_in[1279:1264];
    adder_tree_tier_2_in[655:640] = adder_tree_tier_1_in[1295:1280] + adder_tree_tier_1_in[1311:1296];
    adder_tree_tier_2_in[671:656] = adder_tree_tier_1_in[1327:1312] + adder_tree_tier_1_in[1343:1328];
    adder_tree_tier_2_in[687:672] = adder_tree_tier_1_in[1359:1344] + adder_tree_tier_1_in[1375:1360];
    adder_tree_tier_2_in[703:688] = adder_tree_tier_1_in[1391:1376] + adder_tree_tier_1_in[1407:1392];
    adder_tree_tier_2_in[719:704] = adder_tree_tier_1_in[1423:1408] + adder_tree_tier_1_in[1439:1424];
    adder_tree_tier_2_in[735:720] = adder_tree_tier_1_in[1455:1440] + adder_tree_tier_1_in[1471:1456];
    adder_tree_tier_2_in[751:736] = adder_tree_tier_1_in[1487:1472] + adder_tree_tier_1_in[1503:1488];
    adder_tree_tier_2_in[767:752] = adder_tree_tier_1_in[1519:1504] + adder_tree_tier_1_in[1535:1520];
    adder_tree_tier_2_in[783:768] = adder_tree_tier_1_in[1551:1536] + adder_tree_tier_1_in[1567:1552];
    adder_tree_tier_2_in[799:784] = adder_tree_tier_1_in[1583:1568] + adder_tree_tier_1_in[1599:1584];
    adder_tree_tier_2_in[815:800] = adder_tree_tier_1_in[1615:1600] + adder_tree_tier_1_in[1631:1616];
    adder_tree_tier_2_in[831:816] = adder_tree_tier_1_in[1647:1632] + adder_tree_tier_1_in[1663:1648];
    adder_tree_tier_2_in[847:832] = adder_tree_tier_1_in[1679:1664] + adder_tree_tier_1_in[1695:1680];
    adder_tree_tier_2_in[863:848] = adder_tree_tier_1_in[1711:1696] + adder_tree_tier_1_in[1727:1712];
    adder_tree_tier_2_in[879:864] = adder_tree_tier_1_in[1743:1728] + adder_tree_tier_1_in[1759:1744];
    adder_tree_tier_2_in[895:880] = adder_tree_tier_1_in[1775:1760] + adder_tree_tier_1_in[1791:1776];
    adder_tree_tier_2_in[911:896] = adder_tree_tier_1_in[1807:1792] + adder_tree_tier_1_in[1823:1808];
    adder_tree_tier_2_in[927:912] = adder_tree_tier_1_in[1839:1824] + adder_tree_tier_1_in[1855:1840];
    adder_tree_tier_2_in[943:928] = adder_tree_tier_1_in[1871:1856] + adder_tree_tier_1_in[1887:1872];
    adder_tree_tier_2_in[959:944] = adder_tree_tier_1_in[1903:1888] + adder_tree_tier_1_in[1919:1904];
    adder_tree_tier_2_in[975:960] = adder_tree_tier_1_in[1935:1920] + adder_tree_tier_1_in[1951:1936];
    adder_tree_tier_2_in[991:976] = adder_tree_tier_1_in[1967:1952] + adder_tree_tier_1_in[1983:1968];
    adder_tree_tier_2_in[1007:992] = adder_tree_tier_1_in[1999:1984] + adder_tree_tier_1_in[2015:2000];
    adder_tree_tier_2_in[1023:1008] = adder_tree_tier_1_in[2031:2016] + adder_tree_tier_1_in[2047:2032];
    adder_tree_tier_2_in[1039:1024] = adder_tree_tier_1_in[2063:2048] + adder_tree_tier_1_in[2079:2064];
    adder_tree_tier_2_in[1055:1040] = adder_tree_tier_1_in[2095:2080] + adder_tree_tier_1_in[2111:2096];
    adder_tree_tier_2_in[1071:1056] = adder_tree_tier_1_in[2127:2112] + adder_tree_tier_1_in[2143:2128];
    adder_tree_tier_2_in[1087:1072] = adder_tree_tier_1_in[2159:2144] + adder_tree_tier_1_in[2175:2160];
    adder_tree_tier_2_in[1103:1088] = adder_tree_tier_1_in[2191:2176] + adder_tree_tier_1_in[2207:2192];
    adder_tree_tier_2_in[1119:1104] = adder_tree_tier_1_in[2223:2208] + adder_tree_tier_1_in[2239:2224];
    adder_tree_tier_2_in[1135:1120] = adder_tree_tier_1_in[2255:2240] + adder_tree_tier_1_in[2271:2256];
    adder_tree_tier_2_in[1151:1136] = adder_tree_tier_1_in[2287:2272] + adder_tree_tier_1_in[2303:2288];
    adder_tree_tier_2_in[1167:1152] = adder_tree_tier_1_in[2319:2304] + adder_tree_tier_1_in[2335:2320];
    adder_tree_tier_2_in[1183:1168] = adder_tree_tier_1_in[2351:2336] + adder_tree_tier_1_in[2367:2352];
    adder_tree_tier_2_in[1199:1184] = adder_tree_tier_1_in[2383:2368] + adder_tree_tier_1_in[2399:2384];
    adder_tree_tier_2_in[1215:1200] = adder_tree_tier_1_in[2415:2400] + adder_tree_tier_1_in[2431:2416];
    adder_tree_tier_2_in[1231:1216] = adder_tree_tier_1_in[2447:2432] + adder_tree_tier_1_in[2463:2448];
    adder_tree_tier_2_in[1247:1232] = adder_tree_tier_1_in[2479:2464] + adder_tree_tier_1_in[2495:2480];
    adder_tree_tier_2_in[1263:1248] = adder_tree_tier_1_in[2511:2496] + adder_tree_tier_1_in[2527:2512];
    adder_tree_tier_2_in[1279:1264] = adder_tree_tier_1_in[2543:2528] + adder_tree_tier_1_in[2559:2544];
    adder_tree_tier_2_in[1295:1280] = adder_tree_tier_1_in[2575:2560] + adder_tree_tier_1_in[2591:2576];
    adder_tree_tier_2_in[1311:1296] = adder_tree_tier_1_in[2607:2592] + adder_tree_tier_1_in[2623:2608];
    adder_tree_tier_2_in[1327:1312] = adder_tree_tier_1_in[2639:2624] + adder_tree_tier_1_in[2655:2640];
    adder_tree_tier_2_in[1343:1328] = adder_tree_tier_1_in[2671:2656] + adder_tree_tier_1_in[2687:2672];
    adder_tree_tier_2_in[1359:1344] = adder_tree_tier_1_in[2703:2688] + adder_tree_tier_1_in[2719:2704];
    adder_tree_tier_2_in[1375:1360] = adder_tree_tier_1_in[2735:2720] + adder_tree_tier_1_in[2751:2736];
    adder_tree_tier_2_in[1391:1376] = adder_tree_tier_1_in[2767:2752] + adder_tree_tier_1_in[2783:2768];
    adder_tree_tier_2_in[1407:1392] = adder_tree_tier_1_in[2799:2784] + adder_tree_tier_1_in[2815:2800];
    adder_tree_tier_2_in[1423:1408] = adder_tree_tier_1_in[2831:2816] + adder_tree_tier_1_in[2847:2832];
    adder_tree_tier_2_in[1439:1424] = adder_tree_tier_1_in[2863:2848] + adder_tree_tier_1_in[2879:2864];
    adder_tree_tier_2_in[1455:1440] = adder_tree_tier_1_in[2895:2880] + adder_tree_tier_1_in[2911:2896];
    adder_tree_tier_2_in[1471:1456] = adder_tree_tier_1_in[2927:2912] + adder_tree_tier_1_in[2943:2928];
    adder_tree_tier_2_in[1487:1472] = adder_tree_tier_1_in[2959:2944] + adder_tree_tier_1_in[2975:2960];
    adder_tree_tier_2_in[1503:1488] = adder_tree_tier_1_in[2991:2976] + adder_tree_tier_1_in[3007:2992];
    adder_tree_tier_2_in[1519:1504] = adder_tree_tier_1_in[3023:3008] + adder_tree_tier_1_in[3039:3024];
    adder_tree_tier_2_in[1535:1520] = adder_tree_tier_1_in[3055:3040] + adder_tree_tier_1_in[3071:3056];
    adder_tree_tier_2_in[1551:1536] = adder_tree_tier_1_in[3087:3072] + adder_tree_tier_1_in[3103:3088];
    adder_tree_tier_2_in[1567:1552] = adder_tree_tier_1_in[3119:3104] + adder_tree_tier_1_in[3135:3120];
    adder_tree_tier_2_in[1583:1568] = adder_tree_tier_1_in[3151:3136] + adder_tree_tier_1_in[3167:3152];
    adder_tree_tier_2_in[1599:1584] = adder_tree_tier_1_in[3183:3168] + adder_tree_tier_1_in[3199:3184];
    adder_tree_tier_2_in[1615:1600] = adder_tree_tier_1_in[3215:3200];
    adder_tree_tier_3_in[15:0] = adder_tree_tier_2_in[15:0] + adder_tree_tier_2_in[31:16];
    adder_tree_tier_3_in[31:16] = adder_tree_tier_2_in[47:32] + adder_tree_tier_2_in[63:48];
    adder_tree_tier_3_in[47:32] = adder_tree_tier_2_in[79:64] + adder_tree_tier_2_in[95:80];
    adder_tree_tier_3_in[63:48] = adder_tree_tier_2_in[111:96] + adder_tree_tier_2_in[127:112];
    adder_tree_tier_3_in[79:64] = adder_tree_tier_2_in[143:128] + adder_tree_tier_2_in[159:144];
    adder_tree_tier_3_in[95:80] = adder_tree_tier_2_in[175:160] + adder_tree_tier_2_in[191:176];
    adder_tree_tier_3_in[111:96] = adder_tree_tier_2_in[207:192] + adder_tree_tier_2_in[223:208];
    adder_tree_tier_3_in[127:112] = adder_tree_tier_2_in[239:224] + adder_tree_tier_2_in[255:240];
    adder_tree_tier_3_in[143:128] = adder_tree_tier_2_in[271:256] + adder_tree_tier_2_in[287:272];
    adder_tree_tier_3_in[159:144] = adder_tree_tier_2_in[303:288] + adder_tree_tier_2_in[319:304];
    adder_tree_tier_3_in[175:160] = adder_tree_tier_2_in[335:320] + adder_tree_tier_2_in[351:336];
    adder_tree_tier_3_in[191:176] = adder_tree_tier_2_in[367:352] + adder_tree_tier_2_in[383:368];
    adder_tree_tier_3_in[207:192] = adder_tree_tier_2_in[399:384] + adder_tree_tier_2_in[415:400];
    adder_tree_tier_3_in[223:208] = adder_tree_tier_2_in[431:416] + adder_tree_tier_2_in[447:432];
    adder_tree_tier_3_in[239:224] = adder_tree_tier_2_in[463:448] + adder_tree_tier_2_in[479:464];
    adder_tree_tier_3_in[255:240] = adder_tree_tier_2_in[495:480] + adder_tree_tier_2_in[511:496];
    adder_tree_tier_3_in[271:256] = adder_tree_tier_2_in[527:512] + adder_tree_tier_2_in[543:528];
    adder_tree_tier_3_in[287:272] = adder_tree_tier_2_in[559:544] + adder_tree_tier_2_in[575:560];
    adder_tree_tier_3_in[303:288] = adder_tree_tier_2_in[591:576] + adder_tree_tier_2_in[607:592];
    adder_tree_tier_3_in[319:304] = adder_tree_tier_2_in[623:608] + adder_tree_tier_2_in[639:624];
    adder_tree_tier_3_in[335:320] = adder_tree_tier_2_in[655:640] + adder_tree_tier_2_in[671:656];
    adder_tree_tier_3_in[351:336] = adder_tree_tier_2_in[687:672] + adder_tree_tier_2_in[703:688];
    adder_tree_tier_3_in[367:352] = adder_tree_tier_2_in[719:704] + adder_tree_tier_2_in[735:720];
    adder_tree_tier_3_in[383:368] = adder_tree_tier_2_in[751:736] + adder_tree_tier_2_in[767:752];
    adder_tree_tier_3_in[399:384] = adder_tree_tier_2_in[783:768] + adder_tree_tier_2_in[799:784];
    adder_tree_tier_3_in[415:400] = adder_tree_tier_2_in[815:800] + adder_tree_tier_2_in[831:816];
    adder_tree_tier_3_in[431:416] = adder_tree_tier_2_in[847:832] + adder_tree_tier_2_in[863:848];
    adder_tree_tier_3_in[447:432] = adder_tree_tier_2_in[879:864] + adder_tree_tier_2_in[895:880];
    adder_tree_tier_3_in[463:448] = adder_tree_tier_2_in[911:896] + adder_tree_tier_2_in[927:912];
    adder_tree_tier_3_in[479:464] = adder_tree_tier_2_in[943:928] + adder_tree_tier_2_in[959:944];
    adder_tree_tier_3_in[495:480] = adder_tree_tier_2_in[975:960] + adder_tree_tier_2_in[991:976];
    adder_tree_tier_3_in[511:496] = adder_tree_tier_2_in[1007:992] + adder_tree_tier_2_in[1023:1008];
    adder_tree_tier_3_in[527:512] = adder_tree_tier_2_in[1039:1024] + adder_tree_tier_2_in[1055:1040];
    adder_tree_tier_3_in[543:528] = adder_tree_tier_2_in[1071:1056] + adder_tree_tier_2_in[1087:1072];
    adder_tree_tier_3_in[559:544] = adder_tree_tier_2_in[1103:1088] + adder_tree_tier_2_in[1119:1104];
    adder_tree_tier_3_in[575:560] = adder_tree_tier_2_in[1135:1120] + adder_tree_tier_2_in[1151:1136];
    adder_tree_tier_3_in[591:576] = adder_tree_tier_2_in[1167:1152] + adder_tree_tier_2_in[1183:1168];
    adder_tree_tier_3_in[607:592] = adder_tree_tier_2_in[1199:1184] + adder_tree_tier_2_in[1215:1200];
    adder_tree_tier_3_in[623:608] = adder_tree_tier_2_in[1231:1216] + adder_tree_tier_2_in[1247:1232];
    adder_tree_tier_3_in[639:624] = adder_tree_tier_2_in[1263:1248] + adder_tree_tier_2_in[1279:1264];
    adder_tree_tier_3_in[655:640] = adder_tree_tier_2_in[1295:1280] + adder_tree_tier_2_in[1311:1296];
    adder_tree_tier_3_in[671:656] = adder_tree_tier_2_in[1327:1312] + adder_tree_tier_2_in[1343:1328];
    adder_tree_tier_3_in[687:672] = adder_tree_tier_2_in[1359:1344] + adder_tree_tier_2_in[1375:1360];
    adder_tree_tier_3_in[703:688] = adder_tree_tier_2_in[1391:1376] + adder_tree_tier_2_in[1407:1392];
    adder_tree_tier_3_in[719:704] = adder_tree_tier_2_in[1423:1408] + adder_tree_tier_2_in[1439:1424];
    adder_tree_tier_3_in[735:720] = adder_tree_tier_2_in[1455:1440] + adder_tree_tier_2_in[1471:1456];
    adder_tree_tier_3_in[751:736] = adder_tree_tier_2_in[1487:1472] + adder_tree_tier_2_in[1503:1488];
    adder_tree_tier_3_in[767:752] = adder_tree_tier_2_in[1519:1504] + adder_tree_tier_2_in[1535:1520];
    adder_tree_tier_3_in[783:768] = adder_tree_tier_2_in[1551:1536] + adder_tree_tier_2_in[1567:1552];
    adder_tree_tier_3_in[799:784] = adder_tree_tier_2_in[1583:1568] + adder_tree_tier_2_in[1599:1584];
    adder_tree_tier_3_in[815:800] = adder_tree_tier_2_in[1615:1600];
    adder_tree_tier_4_in[15:0] = adder_tree_tier_3_in[15:0] + adder_tree_tier_3_in[31:16];
    adder_tree_tier_4_in[31:16] = adder_tree_tier_3_in[47:32] + adder_tree_tier_3_in[63:48];
    adder_tree_tier_4_in[47:32] = adder_tree_tier_3_in[79:64] + adder_tree_tier_3_in[95:80];
    adder_tree_tier_4_in[63:48] = adder_tree_tier_3_in[111:96] + adder_tree_tier_3_in[127:112];
    adder_tree_tier_4_in[79:64] = adder_tree_tier_3_in[143:128] + adder_tree_tier_3_in[159:144];
    adder_tree_tier_4_in[95:80] = adder_tree_tier_3_in[175:160] + adder_tree_tier_3_in[191:176];
    adder_tree_tier_4_in[111:96] = adder_tree_tier_3_in[207:192] + adder_tree_tier_3_in[223:208];
    adder_tree_tier_4_in[127:112] = adder_tree_tier_3_in[239:224] + adder_tree_tier_3_in[255:240];
    adder_tree_tier_4_in[143:128] = adder_tree_tier_3_in[271:256] + adder_tree_tier_3_in[287:272];
    adder_tree_tier_4_in[159:144] = adder_tree_tier_3_in[303:288] + adder_tree_tier_3_in[319:304];
    adder_tree_tier_4_in[175:160] = adder_tree_tier_3_in[335:320] + adder_tree_tier_3_in[351:336];
    adder_tree_tier_4_in[191:176] = adder_tree_tier_3_in[367:352] + adder_tree_tier_3_in[383:368];
    adder_tree_tier_4_in[207:192] = adder_tree_tier_3_in[399:384] + adder_tree_tier_3_in[415:400];
    adder_tree_tier_4_in[223:208] = adder_tree_tier_3_in[431:416] + adder_tree_tier_3_in[447:432];
    adder_tree_tier_4_in[239:224] = adder_tree_tier_3_in[463:448] + adder_tree_tier_3_in[479:464];
    adder_tree_tier_4_in[255:240] = adder_tree_tier_3_in[495:480] + adder_tree_tier_3_in[511:496];
    adder_tree_tier_4_in[271:256] = adder_tree_tier_3_in[527:512] + adder_tree_tier_3_in[543:528];
    adder_tree_tier_4_in[287:272] = adder_tree_tier_3_in[559:544] + adder_tree_tier_3_in[575:560];
    adder_tree_tier_4_in[303:288] = adder_tree_tier_3_in[591:576] + adder_tree_tier_3_in[607:592];
    adder_tree_tier_4_in[319:304] = adder_tree_tier_3_in[623:608] + adder_tree_tier_3_in[639:624];
    adder_tree_tier_4_in[335:320] = adder_tree_tier_3_in[655:640] + adder_tree_tier_3_in[671:656];
    adder_tree_tier_4_in[351:336] = adder_tree_tier_3_in[687:672] + adder_tree_tier_3_in[703:688];
    adder_tree_tier_4_in[367:352] = adder_tree_tier_3_in[719:704] + adder_tree_tier_3_in[735:720];
    adder_tree_tier_4_in[383:368] = adder_tree_tier_3_in[751:736] + adder_tree_tier_3_in[767:752];
    adder_tree_tier_4_in[399:384] = adder_tree_tier_3_in[783:768] + adder_tree_tier_3_in[799:784];
    adder_tree_tier_4_in[415:400] = adder_tree_tier_3_in[815:800];
    adder_tree_tier_5_in[15:0] = adder_tree_tier_4_in[15:0] + adder_tree_tier_4_in[31:16];
    adder_tree_tier_5_in[31:16] = adder_tree_tier_4_in[47:32] + adder_tree_tier_4_in[63:48];
    adder_tree_tier_5_in[47:32] = adder_tree_tier_4_in[79:64] + adder_tree_tier_4_in[95:80];
    adder_tree_tier_5_in[63:48] = adder_tree_tier_4_in[111:96] + adder_tree_tier_4_in[127:112];
    adder_tree_tier_5_in[79:64] = adder_tree_tier_4_in[143:128] + adder_tree_tier_4_in[159:144];
    adder_tree_tier_5_in[95:80] = adder_tree_tier_4_in[175:160] + adder_tree_tier_4_in[191:176];
    adder_tree_tier_5_in[111:96] = adder_tree_tier_4_in[207:192] + adder_tree_tier_4_in[223:208];
    adder_tree_tier_5_in[127:112] = adder_tree_tier_4_in[239:224] + adder_tree_tier_4_in[255:240];
    adder_tree_tier_5_in[143:128] = adder_tree_tier_4_in[271:256] + adder_tree_tier_4_in[287:272];
    adder_tree_tier_5_in[159:144] = adder_tree_tier_4_in[303:288] + adder_tree_tier_4_in[319:304];
    adder_tree_tier_5_in[175:160] = adder_tree_tier_4_in[335:320] + adder_tree_tier_4_in[351:336];
    adder_tree_tier_5_in[191:176] = adder_tree_tier_4_in[367:352] + adder_tree_tier_4_in[383:368];
    adder_tree_tier_5_in[207:192] = adder_tree_tier_4_in[399:384] + adder_tree_tier_4_in[415:400];
    adder_tree_tier_6_in[15:0] = adder_tree_tier_5_in[15:0] + adder_tree_tier_5_in[31:16];
    adder_tree_tier_6_in[31:16] = adder_tree_tier_5_in[47:32] + adder_tree_tier_5_in[63:48];
    adder_tree_tier_6_in[47:32] = adder_tree_tier_5_in[79:64] + adder_tree_tier_5_in[95:80];
    adder_tree_tier_6_in[63:48] = adder_tree_tier_5_in[111:96] + adder_tree_tier_5_in[127:112];
    adder_tree_tier_6_in[79:64] = adder_tree_tier_5_in[143:128] + adder_tree_tier_5_in[159:144];
    adder_tree_tier_6_in[95:80] = adder_tree_tier_5_in[175:160] + adder_tree_tier_5_in[191:176];
    adder_tree_tier_6_in[111:96] = adder_tree_tier_5_in[207:192];
    adder_tree_tier_7_in[15:0] = adder_tree_tier_6_in[15:0] + adder_tree_tier_6_in[31:16];
    adder_tree_tier_7_in[31:16] = adder_tree_tier_6_in[47:32] + adder_tree_tier_6_in[63:48];
    adder_tree_tier_7_in[47:32] = adder_tree_tier_6_in[79:64] + adder_tree_tier_6_in[95:80];
    adder_tree_tier_7_in[63:48] = adder_tree_tier_6_in[111:96];
    adder_tree_tier_8_in[15:0] = adder_tree_tier_7_in[15:0] + adder_tree_tier_7_in[31:16];
    adder_tree_tier_8_in[31:16] = adder_tree_tier_7_in[47:32] + adder_tree_tier_7_in[63:48];
    adder_tree_tier_9_in[15:0] = adder_tree_tier_8_in[15:0] + adder_tree_tier_8_in[31:16];
    val_out_buffer = adder_tree_tier_9_in;
  end
  always_ff @(posedge clk or negedge reset) begin
    if (!reset) begin
      history = {(6400){1'b0} };
    end
    else begin
      history = (((history << 16) & {{6384{1'b1}}, {16{1'b0}}}) | cur_val_q);
    end
  end
  always_ff @(posedge clk or negedge reset) begin
    logic [127:0] val_out_buffer_int;
    if (!reset) begin
      val_out_buffer_int = {(143){1'b0} };
    end
    else begin
      val_out_buffer_int = (((val_out_buffer_int << 16) & {{112{1'b1}}, {16{1'b0}}}) | val_out_buffer);
      val_out = val_out_buffer_int[127:112];
    end
  end
endmodule